// Q8.8 Fixed-Point ROM: rom_test_inputs
module rom_test_inputs (
    input [3:0] addr,
    input [10:0] index,
    output reg signed [15:0] data_out
);

    reg signed [15:0] rom [0:9][0:1273];

    initial begin
        rom[0][0] = 16'h0216;
        rom[0][1] = 16'h0162;
        rom[0][2] = 16'h01B8;
        rom[0][3] = 16'h01EB;
        rom[0][4] = 16'h01BF;
        rom[0][5] = 16'h017F;
        rom[0][6] = 16'h014C;
        rom[0][7] = 16'h012F;
        rom[0][8] = 16'h0104;
        rom[0][9] = 16'h00E0;
        rom[0][10] = 16'h00CA;
        rom[0][11] = 16'h00B4;
        rom[0][12] = 16'h00AD;
        rom[0][13] = 16'h00AD;
        rom[0][14] = 16'h009F;
        rom[0][15] = 16'h0098;
        rom[0][16] = 16'h009F;
        rom[0][17] = 16'h00B4;
        rom[0][18] = 16'h00CA;
        rom[0][19] = 16'h00FD;
        rom[0][20] = 16'h0128;
        rom[0][21] = 16'h015A;
        rom[0][22] = 16'h018D;
        rom[0][23] = 16'h0208;
        rom[0][24] = 16'h026D;
        rom[0][25] = 16'h027B;
        rom[0][26] = 16'h0282;
        rom[0][27] = 16'h0291;
        rom[0][28] = 16'h0291;
        rom[0][29] = 16'h0298;
        rom[0][30] = 16'h02A6;
        rom[0][31] = 16'h02B5;
        rom[0][32] = 16'h0000;
        rom[0][33] = 16'h0000;
        rom[0][34] = 16'h0000;
        rom[0][35] = 16'h0000;
        rom[0][36] = 16'h0000;
        rom[0][37] = 16'h0000;
        rom[0][38] = 16'h0000;
        rom[0][39] = 16'h0000;
        rom[0][40] = 16'h0000;
        rom[0][41] = 16'h0000;
        rom[0][42] = 16'h0000;
        rom[0][43] = 16'h0000;
        rom[0][44] = 16'h0000;
        rom[0][45] = 16'h0000;
        rom[0][46] = 16'h0000;
        rom[0][47] = 16'h0000;
        rom[0][48] = 16'h0000;
        rom[0][49] = 16'h0000;
        rom[0][50] = 16'h0000;
        rom[0][51] = 16'h0000;
        rom[0][52] = 16'h0000;
        rom[0][53] = 16'h0000;
        rom[0][54] = 16'h0000;
        rom[0][55] = 16'h0000;
        rom[0][56] = 16'h0000;
        rom[0][57] = 16'h0000;
        rom[0][58] = 16'h0000;
        rom[0][59] = 16'h0000;
        rom[0][60] = 16'h0000;
        rom[0][61] = 16'h0000;
        rom[0][62] = 16'h0000;
        rom[0][63] = 16'h0000;
        rom[0][64] = 16'h0000;
        rom[0][65] = 16'h0000;
        rom[0][66] = 16'h0000;
        rom[0][67] = 16'h0000;
        rom[0][68] = 16'h0000;
        rom[0][69] = 16'h0000;
        rom[0][70] = 16'h0000;
        rom[0][71] = 16'h0000;
        rom[0][72] = 16'h0000;
        rom[0][73] = 16'h0000;
        rom[0][74] = 16'h0000;
        rom[0][75] = 16'h0000;
        rom[0][76] = 16'h0000;
        rom[0][77] = 16'h0000;
        rom[0][78] = 16'h0000;
        rom[0][79] = 16'h0000;
        rom[0][80] = 16'h0000;
        rom[0][81] = 16'h0000;
        rom[0][82] = 16'h0000;
        rom[0][83] = 16'h0000;
        rom[0][84] = 16'h0000;
        rom[0][85] = 16'h0000;
        rom[0][86] = 16'h0000;
        rom[0][87] = 16'h0000;
        rom[0][88] = 16'h0000;
        rom[0][89] = 16'h0000;
        rom[0][90] = 16'h0000;
        rom[0][91] = 16'h0000;
        rom[0][92] = 16'h0000;
        rom[0][93] = 16'h0000;
        rom[0][94] = 16'h0000;
        rom[0][95] = 16'h0000;
        rom[0][96] = 16'h0000;
        rom[0][97] = 16'h0000;
        rom[0][98] = 16'h0177;
        rom[0][99] = 16'h0186;
        rom[0][100] = 16'h00FD;
        rom[0][101] = 16'h009F;
        rom[0][102] = 16'h0065;
        rom[0][103] = 16'h0033;
        rom[0][104] = 16'h000E;
        rom[0][105] = 16'hFFEA;
        rom[0][106] = 16'hFFB8;
        rom[0][107] = 16'hFF94;
        rom[0][108] = 16'hFF7E;
        rom[0][109] = 16'hFF5A;
        rom[0][110] = 16'hFF3D;
        rom[0][111] = 16'hFF5A;
        rom[0][112] = 16'hFF61;
        rom[0][113] = 16'hFF53;
        rom[0][114] = 16'hFF36;
        rom[0][115] = 16'hFF44;
        rom[0][116] = 16'hFF77;
        rom[0][117] = 16'hFF8D;
        rom[0][118] = 16'hFF7E;
        rom[0][119] = 16'hFF7E;
        rom[0][120] = 16'hFFA2;
        rom[0][121] = 16'hFFF9;
        rom[0][122] = 16'h000E;
        rom[0][123] = 16'hFFF9;
        rom[0][124] = 16'h0041;
        rom[0][125] = 16'h00B4;
        rom[0][126] = 16'h0104;
        rom[0][127] = 16'h0121;
        rom[0][128] = 16'h0121;
        rom[0][129] = 16'h013E;
        rom[0][130] = 16'h0000;
        rom[0][131] = 16'h0000;
        rom[0][132] = 16'h0000;
        rom[0][133] = 16'h0000;
        rom[0][134] = 16'h0000;
        rom[0][135] = 16'h0000;
        rom[0][136] = 16'h0000;
        rom[0][137] = 16'h0000;
        rom[0][138] = 16'h0000;
        rom[0][139] = 16'h0000;
        rom[0][140] = 16'h0000;
        rom[0][141] = 16'h0000;
        rom[0][142] = 16'h0000;
        rom[0][143] = 16'h0000;
        rom[0][144] = 16'h0000;
        rom[0][145] = 16'h0000;
        rom[0][146] = 16'h0000;
        rom[0][147] = 16'h0000;
        rom[0][148] = 16'h0000;
        rom[0][149] = 16'h0000;
        rom[0][150] = 16'h0000;
        rom[0][151] = 16'h0000;
        rom[0][152] = 16'h0000;
        rom[0][153] = 16'h0000;
        rom[0][154] = 16'h0000;
        rom[0][155] = 16'h0000;
        rom[0][156] = 16'h0000;
        rom[0][157] = 16'h0000;
        rom[0][158] = 16'h0000;
        rom[0][159] = 16'h0000;
        rom[0][160] = 16'h0000;
        rom[0][161] = 16'h0000;
        rom[0][162] = 16'h0000;
        rom[0][163] = 16'h0000;
        rom[0][164] = 16'h0000;
        rom[0][165] = 16'h0000;
        rom[0][166] = 16'h0000;
        rom[0][167] = 16'h0000;
        rom[0][168] = 16'h0000;
        rom[0][169] = 16'h0000;
        rom[0][170] = 16'h0000;
        rom[0][171] = 16'h0000;
        rom[0][172] = 16'h0000;
        rom[0][173] = 16'h0000;
        rom[0][174] = 16'h0000;
        rom[0][175] = 16'h0000;
        rom[0][176] = 16'h0000;
        rom[0][177] = 16'h0000;
        rom[0][178] = 16'h0000;
        rom[0][179] = 16'h0000;
        rom[0][180] = 16'h0000;
        rom[0][181] = 16'h0000;
        rom[0][182] = 16'h0000;
        rom[0][183] = 16'h0000;
        rom[0][184] = 16'h0000;
        rom[0][185] = 16'h0000;
        rom[0][186] = 16'h0000;
        rom[0][187] = 16'h0000;
        rom[0][188] = 16'h0000;
        rom[0][189] = 16'h0000;
        rom[0][190] = 16'h0000;
        rom[0][191] = 16'h0000;
        rom[0][192] = 16'h0000;
        rom[0][193] = 16'h0000;
        rom[0][194] = 16'h0000;
        rom[0][195] = 16'h0000;
        rom[0][196] = 16'h004F;
        rom[0][197] = 16'h004F;
        rom[0][198] = 16'hFFA2;
        rom[0][199] = 16'hFF94;
        rom[0][200] = 16'hFF9B;
        rom[0][201] = 16'hFF8D;
        rom[0][202] = 16'hFF77;
        rom[0][203] = 16'hFF9B;
        rom[0][204] = 16'hFFA2;
        rom[0][205] = 16'hFFA9;
        rom[0][206] = 16'hFFB1;
        rom[0][207] = 16'hFFA2;
        rom[0][208] = 16'hFF94;
        rom[0][209] = 16'hFFBF;
        rom[0][210] = 16'hFFBF;
        rom[0][211] = 16'hFFC6;
        rom[0][212] = 16'hFFBF;
        rom[0][213] = 16'hFF94;
        rom[0][214] = 16'hFFD5;
        rom[0][215] = 16'hFFD5;
        rom[0][216] = 16'hFFA2;
        rom[0][217] = 16'hFF85;
        rom[0][218] = 16'hFF5A;
        rom[0][219] = 16'hFF20;
        rom[0][220] = 16'hFEFC;
        rom[0][221] = 16'hFEA6;
        rom[0][222] = 16'hFE39;
        rom[0][223] = 16'hFE7A;
        rom[0][224] = 16'hFEC2;
        rom[0][225] = 16'hFF0B;
        rom[0][226] = 16'hFEEE;
        rom[0][227] = 16'hFE97;
        rom[0][228] = 16'h0000;
        rom[0][229] = 16'h0000;
        rom[0][230] = 16'h0000;
        rom[0][231] = 16'h0000;
        rom[0][232] = 16'h0000;
        rom[0][233] = 16'h0000;
        rom[0][234] = 16'h0000;
        rom[0][235] = 16'h0000;
        rom[0][236] = 16'h0000;
        rom[0][237] = 16'h0000;
        rom[0][238] = 16'h0000;
        rom[0][239] = 16'h0000;
        rom[0][240] = 16'h0000;
        rom[0][241] = 16'h0000;
        rom[0][242] = 16'h0000;
        rom[0][243] = 16'h0000;
        rom[0][244] = 16'h0000;
        rom[0][245] = 16'h0000;
        rom[0][246] = 16'h0000;
        rom[0][247] = 16'h0000;
        rom[0][248] = 16'h0000;
        rom[0][249] = 16'h0000;
        rom[0][250] = 16'h0000;
        rom[0][251] = 16'h0000;
        rom[0][252] = 16'h0000;
        rom[0][253] = 16'h0000;
        rom[0][254] = 16'h0000;
        rom[0][255] = 16'h0000;
        rom[0][256] = 16'h0000;
        rom[0][257] = 16'h0000;
        rom[0][258] = 16'h0000;
        rom[0][259] = 16'h0000;
        rom[0][260] = 16'h0000;
        rom[0][261] = 16'h0000;
        rom[0][262] = 16'h0000;
        rom[0][263] = 16'h0000;
        rom[0][264] = 16'h0000;
        rom[0][265] = 16'h0000;
        rom[0][266] = 16'h0000;
        rom[0][267] = 16'h0000;
        rom[0][268] = 16'h0000;
        rom[0][269] = 16'h0000;
        rom[0][270] = 16'h0000;
        rom[0][271] = 16'h0000;
        rom[0][272] = 16'h0000;
        rom[0][273] = 16'h0000;
        rom[0][274] = 16'h0000;
        rom[0][275] = 16'h0000;
        rom[0][276] = 16'h0000;
        rom[0][277] = 16'h0000;
        rom[0][278] = 16'h0000;
        rom[0][279] = 16'h0000;
        rom[0][280] = 16'h0000;
        rom[0][281] = 16'h0000;
        rom[0][282] = 16'h0000;
        rom[0][283] = 16'h0000;
        rom[0][284] = 16'h0000;
        rom[0][285] = 16'h0000;
        rom[0][286] = 16'h0000;
        rom[0][287] = 16'h0000;
        rom[0][288] = 16'h0000;
        rom[0][289] = 16'h0000;
        rom[0][290] = 16'h0000;
        rom[0][291] = 16'h0000;
        rom[0][292] = 16'h0000;
        rom[0][293] = 16'h0000;
        rom[0][294] = 16'hFF53;
        rom[0][295] = 16'hFEFC;
        rom[0][296] = 16'hFE81;
        rom[0][297] = 16'hFE73;
        rom[0][298] = 16'hFE9E;
        rom[0][299] = 16'hFE97;
        rom[0][300] = 16'hFE9E;
        rom[0][301] = 16'hFE81;
        rom[0][302] = 16'hFE7A;
        rom[0][303] = 16'hFE65;
        rom[0][304] = 16'hFE7A;
        rom[0][305] = 16'hFE73;
        rom[0][306] = 16'hFE9E;
        rom[0][307] = 16'hFEFC;
        rom[0][308] = 16'hFEE7;
        rom[0][309] = 16'hFEBB;
        rom[0][310] = 16'hFEAD;
        rom[0][311] = 16'hFEAD;
        rom[0][312] = 16'hFF3D;
        rom[0][313] = 16'h0000;
        rom[0][314] = 16'h0048;
        rom[0][315] = 16'h0041;
        rom[0][316] = 16'h000E;
        rom[0][317] = 16'h001D;
        rom[0][318] = 16'hFFF9;
        rom[0][319] = 16'hFF9B;
        rom[0][320] = 16'hFEFC;
        rom[0][321] = 16'hFEB4;
        rom[0][322] = 16'hFE81;
        rom[0][323] = 16'hFE81;
        rom[0][324] = 16'hFE2B;
        rom[0][325] = 16'hFDEA;
        rom[0][326] = 16'h0000;
        rom[0][327] = 16'h0000;
        rom[0][328] = 16'h0000;
        rom[0][329] = 16'h0000;
        rom[0][330] = 16'h0000;
        rom[0][331] = 16'h0000;
        rom[0][332] = 16'h0000;
        rom[0][333] = 16'h0000;
        rom[0][334] = 16'h0000;
        rom[0][335] = 16'h0000;
        rom[0][336] = 16'h0000;
        rom[0][337] = 16'h0000;
        rom[0][338] = 16'h0000;
        rom[0][339] = 16'h0000;
        rom[0][340] = 16'h0000;
        rom[0][341] = 16'h0000;
        rom[0][342] = 16'h0000;
        rom[0][343] = 16'h0000;
        rom[0][344] = 16'h0000;
        rom[0][345] = 16'h0000;
        rom[0][346] = 16'h0000;
        rom[0][347] = 16'h0000;
        rom[0][348] = 16'h0000;
        rom[0][349] = 16'h0000;
        rom[0][350] = 16'h0000;
        rom[0][351] = 16'h0000;
        rom[0][352] = 16'h0000;
        rom[0][353] = 16'h0000;
        rom[0][354] = 16'h0000;
        rom[0][355] = 16'h0000;
        rom[0][356] = 16'h0000;
        rom[0][357] = 16'h0000;
        rom[0][358] = 16'h0000;
        rom[0][359] = 16'h0000;
        rom[0][360] = 16'h0000;
        rom[0][361] = 16'h0000;
        rom[0][362] = 16'h0000;
        rom[0][363] = 16'h0000;
        rom[0][364] = 16'h0000;
        rom[0][365] = 16'h0000;
        rom[0][366] = 16'h0000;
        rom[0][367] = 16'h0000;
        rom[0][368] = 16'h0000;
        rom[0][369] = 16'h0000;
        rom[0][370] = 16'h0000;
        rom[0][371] = 16'h0000;
        rom[0][372] = 16'h0000;
        rom[0][373] = 16'h0000;
        rom[0][374] = 16'h0000;
        rom[0][375] = 16'h0000;
        rom[0][376] = 16'h0000;
        rom[0][377] = 16'h0000;
        rom[0][378] = 16'h0000;
        rom[0][379] = 16'h0000;
        rom[0][380] = 16'h0000;
        rom[0][381] = 16'h0000;
        rom[0][382] = 16'h0000;
        rom[0][383] = 16'h0000;
        rom[0][384] = 16'h0000;
        rom[0][385] = 16'h0000;
        rom[0][386] = 16'h0000;
        rom[0][387] = 16'h0000;
        rom[0][388] = 16'h0000;
        rom[0][389] = 16'h0000;
        rom[0][390] = 16'h0000;
        rom[0][391] = 16'h0000;
        rom[0][392] = 16'hFE81;
        rom[0][393] = 16'hFE24;
        rom[0][394] = 16'hFD7E;
        rom[0][395] = 16'hFE07;
        rom[0][396] = 16'hFE1C;
        rom[0][397] = 16'hFE24;
        rom[0][398] = 16'hFE90;
        rom[0][399] = 16'hFED1;
        rom[0][400] = 16'hFED1;
        rom[0][401] = 16'hFE81;
        rom[0][402] = 16'hFEBB;
        rom[0][403] = 16'hFED1;
        rom[0][404] = 16'hFEE7;
        rom[0][405] = 16'hFF5A;
        rom[0][406] = 16'hFF7E;
        rom[0][407] = 16'hFF3D;
        rom[0][408] = 16'hFF27;
        rom[0][409] = 16'hFF61;
        rom[0][410] = 16'hFFEA;
        rom[0][411] = 16'h0090;
        rom[0][412] = 16'h00CA;
        rom[0][413] = 16'h0089;
        rom[0][414] = 16'h006C;
        rom[0][415] = 16'hFFE3;
        rom[0][416] = 16'hFF61;
        rom[0][417] = 16'hFEEE;
        rom[0][418] = 16'hFE48;
        rom[0][419] = 16'hFD6F;
        rom[0][420] = 16'hFCFC;
        rom[0][421] = 16'hFD11;
        rom[0][422] = 16'hFD11;
        rom[0][423] = 16'hFD85;
        rom[0][424] = 16'h0000;
        rom[0][425] = 16'h0000;
        rom[0][426] = 16'h0000;
        rom[0][427] = 16'h0000;
        rom[0][428] = 16'h0000;
        rom[0][429] = 16'h0000;
        rom[0][430] = 16'h0000;
        rom[0][431] = 16'h0000;
        rom[0][432] = 16'h0000;
        rom[0][433] = 16'h0000;
        rom[0][434] = 16'h0000;
        rom[0][435] = 16'h0000;
        rom[0][436] = 16'h0000;
        rom[0][437] = 16'h0000;
        rom[0][438] = 16'h0000;
        rom[0][439] = 16'h0000;
        rom[0][440] = 16'h0000;
        rom[0][441] = 16'h0000;
        rom[0][442] = 16'h0000;
        rom[0][443] = 16'h0000;
        rom[0][444] = 16'h0000;
        rom[0][445] = 16'h0000;
        rom[0][446] = 16'h0000;
        rom[0][447] = 16'h0000;
        rom[0][448] = 16'h0000;
        rom[0][449] = 16'h0000;
        rom[0][450] = 16'h0000;
        rom[0][451] = 16'h0000;
        rom[0][452] = 16'h0000;
        rom[0][453] = 16'h0000;
        rom[0][454] = 16'h0000;
        rom[0][455] = 16'h0000;
        rom[0][456] = 16'h0000;
        rom[0][457] = 16'h0000;
        rom[0][458] = 16'h0000;
        rom[0][459] = 16'h0000;
        rom[0][460] = 16'h0000;
        rom[0][461] = 16'h0000;
        rom[0][462] = 16'h0000;
        rom[0][463] = 16'h0000;
        rom[0][464] = 16'h0000;
        rom[0][465] = 16'h0000;
        rom[0][466] = 16'h0000;
        rom[0][467] = 16'h0000;
        rom[0][468] = 16'h0000;
        rom[0][469] = 16'h0000;
        rom[0][470] = 16'h0000;
        rom[0][471] = 16'h0000;
        rom[0][472] = 16'h0000;
        rom[0][473] = 16'h0000;
        rom[0][474] = 16'h0000;
        rom[0][475] = 16'h0000;
        rom[0][476] = 16'h0000;
        rom[0][477] = 16'h0000;
        rom[0][478] = 16'h0000;
        rom[0][479] = 16'h0000;
        rom[0][480] = 16'h0000;
        rom[0][481] = 16'h0000;
        rom[0][482] = 16'h0000;
        rom[0][483] = 16'h0000;
        rom[0][484] = 16'h0000;
        rom[0][485] = 16'h0000;
        rom[0][486] = 16'h0000;
        rom[0][487] = 16'h0000;
        rom[0][488] = 16'h0000;
        rom[0][489] = 16'h0000;
        rom[0][490] = 16'hFE00;
        rom[0][491] = 16'hFDD4;
        rom[0][492] = 16'hFD11;
        rom[0][493] = 16'hFD61;
        rom[0][494] = 16'hFD93;
        rom[0][495] = 16'hFD7E;
        rom[0][496] = 16'hFDD4;
        rom[0][497] = 16'hFE48;
        rom[0][498] = 16'hFE2B;
        rom[0][499] = 16'hFE00;
        rom[0][500] = 16'hFDDB;
        rom[0][501] = 16'hFDF8;
        rom[0][502] = 16'hFE15;
        rom[0][503] = 16'hFE89;
        rom[0][504] = 16'hFED1;
        rom[0][505] = 16'hFE97;
        rom[0][506] = 16'hFE65;
        rom[0][507] = 16'hFE56;
        rom[0][508] = 16'hFE89;
        rom[0][509] = 16'hFE41;
        rom[0][510] = 16'hFE15;
        rom[0][511] = 16'hFDE3;
        rom[0][512] = 16'hFE07;
        rom[0][513] = 16'hFD4B;
        rom[0][514] = 16'hFD44;
        rom[0][515] = 16'hFDA9;
        rom[0][516] = 16'hFDB0;
        rom[0][517] = 16'hFD27;
        rom[0][518] = 16'h037F;
        rom[0][519] = 16'hFC64;
        rom[0][520] = 16'hFCE6;
        rom[0][521] = 16'hFD44;
        rom[0][522] = 16'h0000;
        rom[0][523] = 16'h0000;
        rom[0][524] = 16'h0000;
        rom[0][525] = 16'h0000;
        rom[0][526] = 16'h0000;
        rom[0][527] = 16'h0000;
        rom[0][528] = 16'h0000;
        rom[0][529] = 16'h0000;
        rom[0][530] = 16'h0000;
        rom[0][531] = 16'h0000;
        rom[0][532] = 16'h0000;
        rom[0][533] = 16'h0000;
        rom[0][534] = 16'h0000;
        rom[0][535] = 16'h0000;
        rom[0][536] = 16'h0000;
        rom[0][537] = 16'h0000;
        rom[0][538] = 16'h0000;
        rom[0][539] = 16'h0000;
        rom[0][540] = 16'h0000;
        rom[0][541] = 16'h0000;
        rom[0][542] = 16'h0000;
        rom[0][543] = 16'h0000;
        rom[0][544] = 16'h0000;
        rom[0][545] = 16'h0000;
        rom[0][546] = 16'h0000;
        rom[0][547] = 16'h0000;
        rom[0][548] = 16'h0000;
        rom[0][549] = 16'h0000;
        rom[0][550] = 16'h0000;
        rom[0][551] = 16'h0000;
        rom[0][552] = 16'h0000;
        rom[0][553] = 16'h0000;
        rom[0][554] = 16'h0000;
        rom[0][555] = 16'h0000;
        rom[0][556] = 16'h0000;
        rom[0][557] = 16'h0000;
        rom[0][558] = 16'h0000;
        rom[0][559] = 16'h0000;
        rom[0][560] = 16'h0000;
        rom[0][561] = 16'h0000;
        rom[0][562] = 16'h0000;
        rom[0][563] = 16'h0000;
        rom[0][564] = 16'h0000;
        rom[0][565] = 16'h0000;
        rom[0][566] = 16'h0000;
        rom[0][567] = 16'h0000;
        rom[0][568] = 16'h0000;
        rom[0][569] = 16'h0000;
        rom[0][570] = 16'h0000;
        rom[0][571] = 16'h0000;
        rom[0][572] = 16'h0000;
        rom[0][573] = 16'h0000;
        rom[0][574] = 16'h0000;
        rom[0][575] = 16'h0000;
        rom[0][576] = 16'h0000;
        rom[0][577] = 16'h0000;
        rom[0][578] = 16'h0000;
        rom[0][579] = 16'h0000;
        rom[0][580] = 16'h0000;
        rom[0][581] = 16'h0000;
        rom[0][582] = 16'h0000;
        rom[0][583] = 16'h0000;
        rom[0][584] = 16'h0000;
        rom[0][585] = 16'h0000;
        rom[0][586] = 16'h0000;
        rom[0][587] = 16'h0000;
        rom[0][588] = 16'hFE73;
        rom[0][589] = 16'hFE73;
        rom[0][590] = 16'hFD85;
        rom[0][591] = 16'hFD9B;
        rom[0][592] = 16'hFDDB;
        rom[0][593] = 16'hFDF8;
        rom[0][594] = 16'hFE00;
        rom[0][595] = 16'hFE5D;
        rom[0][596] = 16'hFE56;
        rom[0][597] = 16'hFE65;
        rom[0][598] = 16'hFE41;
        rom[0][599] = 16'hFE24;
        rom[0][600] = 16'hFE81;
        rom[0][601] = 16'hFEDF;
        rom[0][602] = 16'hFF20;
        rom[0][603] = 16'hFEF5;
        rom[0][604] = 16'hFEC2;
        rom[0][605] = 16'hFEFC;
        rom[0][606] = 16'hFEDF;
        rom[0][607] = 16'hFDD4;
        rom[0][608] = 16'hFD68;
        rom[0][609] = 16'hFD8C;
        rom[0][610] = 16'hFDE3;
        rom[0][611] = 16'hFD93;
        rom[0][612] = 16'hFDA2;
        rom[0][613] = 16'hFD9B;
        rom[0][614] = 16'hFD5A;
        rom[0][615] = 16'hFD2E;
        rom[0][616] = 16'hFCFC;
        rom[0][617] = 16'hFCFC;
        rom[0][618] = 16'hFCF5;
        rom[0][619] = 16'hFCFC;
        rom[0][620] = 16'h0000;
        rom[0][621] = 16'h0000;
        rom[0][622] = 16'h0000;
        rom[0][623] = 16'h0000;
        rom[0][624] = 16'h0000;
        rom[0][625] = 16'h0000;
        rom[0][626] = 16'h0000;
        rom[0][627] = 16'h0000;
        rom[0][628] = 16'h0000;
        rom[0][629] = 16'h0000;
        rom[0][630] = 16'h0000;
        rom[0][631] = 16'h0000;
        rom[0][632] = 16'h0000;
        rom[0][633] = 16'h0000;
        rom[0][634] = 16'h0000;
        rom[0][635] = 16'h0000;
        rom[0][636] = 16'h0000;
        rom[0][637] = 16'h0000;
        rom[0][638] = 16'h0000;
        rom[0][639] = 16'h0000;
        rom[0][640] = 16'h0000;
        rom[0][641] = 16'h0000;
        rom[0][642] = 16'h0000;
        rom[0][643] = 16'h0000;
        rom[0][644] = 16'h0000;
        rom[0][645] = 16'h0000;
        rom[0][646] = 16'h0000;
        rom[0][647] = 16'h0000;
        rom[0][648] = 16'h0000;
        rom[0][649] = 16'h0000;
        rom[0][650] = 16'h0000;
        rom[0][651] = 16'h0000;
        rom[0][652] = 16'h0000;
        rom[0][653] = 16'h0000;
        rom[0][654] = 16'h0000;
        rom[0][655] = 16'h0000;
        rom[0][656] = 16'h0000;
        rom[0][657] = 16'h0000;
        rom[0][658] = 16'h0000;
        rom[0][659] = 16'h0000;
        rom[0][660] = 16'h0000;
        rom[0][661] = 16'h0000;
        rom[0][662] = 16'h0000;
        rom[0][663] = 16'h0000;
        rom[0][664] = 16'h0000;
        rom[0][665] = 16'h0000;
        rom[0][666] = 16'h0000;
        rom[0][667] = 16'h0000;
        rom[0][668] = 16'h0000;
        rom[0][669] = 16'h0000;
        rom[0][670] = 16'h0000;
        rom[0][671] = 16'h0000;
        rom[0][672] = 16'h0000;
        rom[0][673] = 16'h0000;
        rom[0][674] = 16'h0000;
        rom[0][675] = 16'h0000;
        rom[0][676] = 16'h0000;
        rom[0][677] = 16'h0000;
        rom[0][678] = 16'h0000;
        rom[0][679] = 16'h0000;
        rom[0][680] = 16'h0000;
        rom[0][681] = 16'h0000;
        rom[0][682] = 16'h0000;
        rom[0][683] = 16'h0000;
        rom[0][684] = 16'h0000;
        rom[0][685] = 16'h0000;
        rom[0][686] = 16'hFE24;
        rom[0][687] = 16'hFE2B;
        rom[0][688] = 16'hFE73;
        rom[0][689] = 16'hFEAD;
        rom[0][690] = 16'hFE81;
        rom[0][691] = 16'hFE7A;
        rom[0][692] = 16'hFED1;
        rom[0][693] = 16'hFED1;
        rom[0][694] = 16'hFE89;
        rom[0][695] = 16'hFE56;
        rom[0][696] = 16'hFE97;
        rom[0][697] = 16'hFEAD;
        rom[0][698] = 16'hFF0B;
        rom[0][699] = 16'hFF3D;
        rom[0][700] = 16'hFF77;
        rom[0][701] = 16'hFF68;
        rom[0][702] = 16'hFF2F;
        rom[0][703] = 16'hFF3D;
        rom[0][704] = 16'hFF4C;
        rom[0][705] = 16'hFF3D;
        rom[0][706] = 16'hFF0B;
        rom[0][707] = 16'hFFD5;
        rom[0][708] = 16'h001D;
        rom[0][709] = 16'hFF03;
        rom[0][710] = 16'hFE81;
        rom[0][711] = 16'hFEE7;
        rom[0][712] = 16'hFF68;
        rom[0][713] = 16'hFF68;
        rom[0][714] = 16'hFE56;
        rom[0][715] = 16'hFDA2;
        rom[0][716] = 16'hFD93;
        rom[0][717] = 16'hFD35;
        rom[0][718] = 16'h0000;
        rom[0][719] = 16'h0000;
        rom[0][720] = 16'h0000;
        rom[0][721] = 16'h0000;
        rom[0][722] = 16'h0000;
        rom[0][723] = 16'h0000;
        rom[0][724] = 16'h0000;
        rom[0][725] = 16'h0000;
        rom[0][726] = 16'h0000;
        rom[0][727] = 16'h0000;
        rom[0][728] = 16'h0000;
        rom[0][729] = 16'h0000;
        rom[0][730] = 16'h0000;
        rom[0][731] = 16'h0000;
        rom[0][732] = 16'h0000;
        rom[0][733] = 16'h0000;
        rom[0][734] = 16'h0000;
        rom[0][735] = 16'h0000;
        rom[0][736] = 16'h0000;
        rom[0][737] = 16'h0000;
        rom[0][738] = 16'h0000;
        rom[0][739] = 16'h0000;
        rom[0][740] = 16'h0000;
        rom[0][741] = 16'h0000;
        rom[0][742] = 16'h0000;
        rom[0][743] = 16'h0000;
        rom[0][744] = 16'h0000;
        rom[0][745] = 16'h0000;
        rom[0][746] = 16'h0000;
        rom[0][747] = 16'h0000;
        rom[0][748] = 16'h0000;
        rom[0][749] = 16'h0000;
        rom[0][750] = 16'h0000;
        rom[0][751] = 16'h0000;
        rom[0][752] = 16'h0000;
        rom[0][753] = 16'h0000;
        rom[0][754] = 16'h0000;
        rom[0][755] = 16'h0000;
        rom[0][756] = 16'h0000;
        rom[0][757] = 16'h0000;
        rom[0][758] = 16'h0000;
        rom[0][759] = 16'h0000;
        rom[0][760] = 16'h0000;
        rom[0][761] = 16'h0000;
        rom[0][762] = 16'h0000;
        rom[0][763] = 16'h0000;
        rom[0][764] = 16'h0000;
        rom[0][765] = 16'h0000;
        rom[0][766] = 16'h0000;
        rom[0][767] = 16'h0000;
        rom[0][768] = 16'h0000;
        rom[0][769] = 16'h0000;
        rom[0][770] = 16'h0000;
        rom[0][771] = 16'h0000;
        rom[0][772] = 16'h0000;
        rom[0][773] = 16'h0000;
        rom[0][774] = 16'h0000;
        rom[0][775] = 16'h0000;
        rom[0][776] = 16'h0000;
        rom[0][777] = 16'h0000;
        rom[0][778] = 16'h0000;
        rom[0][779] = 16'h0000;
        rom[0][780] = 16'h0000;
        rom[0][781] = 16'h0000;
        rom[0][782] = 16'h0000;
        rom[0][783] = 16'h0000;
        rom[0][784] = 16'hFE15;
        rom[0][785] = 16'hFE56;
        rom[0][786] = 16'hFE00;
        rom[0][787] = 16'hFE00;
        rom[0][788] = 16'hFDCD;
        rom[0][789] = 16'hFE48;
        rom[0][790] = 16'hFEAD;
        rom[0][791] = 16'hFE6C;
        rom[0][792] = 16'hFE41;
        rom[0][793] = 16'hFE41;
        rom[0][794] = 16'hFE97;
        rom[0][795] = 16'hFE5D;
        rom[0][796] = 16'hFE65;
        rom[0][797] = 16'hFE39;
        rom[0][798] = 16'hFE07;
        rom[0][799] = 16'hFE65;
        rom[0][800] = 16'hFE90;
        rom[0][801] = 16'hFEC2;
        rom[0][802] = 16'hFE9E;
        rom[0][803] = 16'hFE0E;
        rom[0][804] = 16'hFD52;
        rom[0][805] = 16'hFD19;
        rom[0][806] = 16'hFD20;
        rom[0][807] = 16'hFEE7;
        rom[0][808] = 16'hFFB8;
        rom[0][809] = 16'hFF77;
        rom[0][810] = 16'hFEAD;
        rom[0][811] = 16'hFDB7;
        rom[0][812] = 16'hFD11;
        rom[0][813] = 16'hFC88;
        rom[0][814] = 16'hFCDF;
        rom[0][815] = 16'hFD93;
        rom[0][816] = 16'h0000;
        rom[0][817] = 16'h0000;
        rom[0][818] = 16'h0000;
        rom[0][819] = 16'h0000;
        rom[0][820] = 16'h0000;
        rom[0][821] = 16'h0000;
        rom[0][822] = 16'h0000;
        rom[0][823] = 16'h0000;
        rom[0][824] = 16'h0000;
        rom[0][825] = 16'h0000;
        rom[0][826] = 16'h0000;
        rom[0][827] = 16'h0000;
        rom[0][828] = 16'h0000;
        rom[0][829] = 16'h0000;
        rom[0][830] = 16'h0000;
        rom[0][831] = 16'h0000;
        rom[0][832] = 16'h0000;
        rom[0][833] = 16'h0000;
        rom[0][834] = 16'h0000;
        rom[0][835] = 16'h0000;
        rom[0][836] = 16'h0000;
        rom[0][837] = 16'h0000;
        rom[0][838] = 16'h0000;
        rom[0][839] = 16'h0000;
        rom[0][840] = 16'h0000;
        rom[0][841] = 16'h0000;
        rom[0][842] = 16'h0000;
        rom[0][843] = 16'h0000;
        rom[0][844] = 16'h0000;
        rom[0][845] = 16'h0000;
        rom[0][846] = 16'h0000;
        rom[0][847] = 16'h0000;
        rom[0][848] = 16'h0000;
        rom[0][849] = 16'h0000;
        rom[0][850] = 16'h0000;
        rom[0][851] = 16'h0000;
        rom[0][852] = 16'h0000;
        rom[0][853] = 16'h0000;
        rom[0][854] = 16'h0000;
        rom[0][855] = 16'h0000;
        rom[0][856] = 16'h0000;
        rom[0][857] = 16'h0000;
        rom[0][858] = 16'h0000;
        rom[0][859] = 16'h0000;
        rom[0][860] = 16'h0000;
        rom[0][861] = 16'h0000;
        rom[0][862] = 16'h0000;
        rom[0][863] = 16'h0000;
        rom[0][864] = 16'h0000;
        rom[0][865] = 16'h0000;
        rom[0][866] = 16'h0000;
        rom[0][867] = 16'h0000;
        rom[0][868] = 16'h0000;
        rom[0][869] = 16'h0000;
        rom[0][870] = 16'h0000;
        rom[0][871] = 16'h0000;
        rom[0][872] = 16'h0000;
        rom[0][873] = 16'h0000;
        rom[0][874] = 16'h0000;
        rom[0][875] = 16'h0000;
        rom[0][876] = 16'h0000;
        rom[0][877] = 16'h0000;
        rom[0][878] = 16'h0000;
        rom[0][879] = 16'h0000;
        rom[0][880] = 16'h0000;
        rom[0][881] = 16'h0000;
        rom[0][882] = 16'hFE39;
        rom[0][883] = 16'hFE65;
        rom[0][884] = 16'hFE2B;
        rom[0][885] = 16'hFE81;
        rom[0][886] = 16'hFE56;
        rom[0][887] = 16'hFE7A;
        rom[0][888] = 16'hFF27;
        rom[0][889] = 16'hFF12;
        rom[0][890] = 16'hFEBB;
        rom[0][891] = 16'hFE97;
        rom[0][892] = 16'hFE7A;
        rom[0][893] = 16'hFEB4;
        rom[0][894] = 16'hFF53;
        rom[0][895] = 16'hFF3D;
        rom[0][896] = 16'hFEEE;
        rom[0][897] = 16'hFF0B;
        rom[0][898] = 16'hFF36;
        rom[0][899] = 16'hFF61;
        rom[0][900] = 16'hFF19;
        rom[0][901] = 16'hFF0B;
        rom[0][902] = 16'hFEFC;
        rom[0][903] = 16'hFF03;
        rom[0][904] = 16'hFEFC;
        rom[0][905] = 16'h00B4;
        rom[0][906] = 16'h014C;
        rom[0][907] = 16'h0169;
        rom[0][908] = 16'h0119;
        rom[0][909] = 16'h00BC;
        rom[0][910] = 16'h00A6;
        rom[0][911] = 16'h00CA;
        rom[0][912] = 16'h005E;
        rom[0][913] = 16'h007B;
        rom[0][914] = 16'h0000;
        rom[0][915] = 16'h0000;
        rom[0][916] = 16'h0000;
        rom[0][917] = 16'h0000;
        rom[0][918] = 16'h0000;
        rom[0][919] = 16'h0000;
        rom[0][920] = 16'h0000;
        rom[0][921] = 16'h0000;
        rom[0][922] = 16'h0000;
        rom[0][923] = 16'h0000;
        rom[0][924] = 16'h0000;
        rom[0][925] = 16'h0000;
        rom[0][926] = 16'h0000;
        rom[0][927] = 16'h0000;
        rom[0][928] = 16'h0000;
        rom[0][929] = 16'h0000;
        rom[0][930] = 16'h0000;
        rom[0][931] = 16'h0000;
        rom[0][932] = 16'h0000;
        rom[0][933] = 16'h0000;
        rom[0][934] = 16'h0000;
        rom[0][935] = 16'h0000;
        rom[0][936] = 16'h0000;
        rom[0][937] = 16'h0000;
        rom[0][938] = 16'h0000;
        rom[0][939] = 16'h0000;
        rom[0][940] = 16'h0000;
        rom[0][941] = 16'h0000;
        rom[0][942] = 16'h0000;
        rom[0][943] = 16'h0000;
        rom[0][944] = 16'h0000;
        rom[0][945] = 16'h0000;
        rom[0][946] = 16'h0000;
        rom[0][947] = 16'h0000;
        rom[0][948] = 16'h0000;
        rom[0][949] = 16'h0000;
        rom[0][950] = 16'h0000;
        rom[0][951] = 16'h0000;
        rom[0][952] = 16'h0000;
        rom[0][953] = 16'h0000;
        rom[0][954] = 16'h0000;
        rom[0][955] = 16'h0000;
        rom[0][956] = 16'h0000;
        rom[0][957] = 16'h0000;
        rom[0][958] = 16'h0000;
        rom[0][959] = 16'h0000;
        rom[0][960] = 16'h0000;
        rom[0][961] = 16'h0000;
        rom[0][962] = 16'h0000;
        rom[0][963] = 16'h0000;
        rom[0][964] = 16'h0000;
        rom[0][965] = 16'h0000;
        rom[0][966] = 16'h0000;
        rom[0][967] = 16'h0000;
        rom[0][968] = 16'h0000;
        rom[0][969] = 16'h0000;
        rom[0][970] = 16'h0000;
        rom[0][971] = 16'h0000;
        rom[0][972] = 16'h0000;
        rom[0][973] = 16'h0000;
        rom[0][974] = 16'h0000;
        rom[0][975] = 16'h0000;
        rom[0][976] = 16'h0000;
        rom[0][977] = 16'h0000;
        rom[0][978] = 16'h0000;
        rom[0][979] = 16'h0000;
        rom[0][980] = 16'hFF85;
        rom[0][981] = 16'hFF68;
        rom[0][982] = 16'hFE39;
        rom[0][983] = 16'hFE4F;
        rom[0][984] = 16'hFEC2;
        rom[0][985] = 16'hFEC2;
        rom[0][986] = 16'hFEEE;
        rom[0][987] = 16'hFF61;
        rom[0][988] = 16'hFF7E;
        rom[0][989] = 16'hFF0B;
        rom[0][990] = 16'hFEDF;
        rom[0][991] = 16'hFF19;
        rom[0][992] = 16'hFFE3;
        rom[0][993] = 16'h0000;
        rom[0][994] = 16'hFF53;
        rom[0][995] = 16'hFF8D;
        rom[0][996] = 16'hFFE3;
        rom[0][997] = 16'hFFEA;
        rom[0][998] = 16'hFFF9;
        rom[0][999] = 16'h001D;
        rom[0][1000] = 16'h001D;
        rom[0][1001] = 16'hFFDC;
        rom[0][1002] = 16'h0024;
        rom[0][1003] = 16'h007B;
        rom[0][1004] = 16'h0082;
        rom[0][1005] = 16'h00CA;
        rom[0][1006] = 16'h0112;
        rom[0][1007] = 16'h0104;
        rom[0][1008] = 16'h00D1;
        rom[0][1009] = 16'h0073;
        rom[0][1010] = 16'hFF85;
        rom[0][1011] = 16'hFF27;
        rom[0][1012] = 16'h0000;
        rom[0][1013] = 16'h0000;
        rom[0][1014] = 16'h0000;
        rom[0][1015] = 16'h0000;
        rom[0][1016] = 16'h0000;
        rom[0][1017] = 16'h0000;
        rom[0][1018] = 16'h0000;
        rom[0][1019] = 16'h0000;
        rom[0][1020] = 16'h0000;
        rom[0][1021] = 16'h0000;
        rom[0][1022] = 16'h0000;
        rom[0][1023] = 16'h0000;
        rom[0][1024] = 16'h0000;
        rom[0][1025] = 16'h0000;
        rom[0][1026] = 16'h0000;
        rom[0][1027] = 16'h0000;
        rom[0][1028] = 16'h0000;
        rom[0][1029] = 16'h0000;
        rom[0][1030] = 16'h0000;
        rom[0][1031] = 16'h0000;
        rom[0][1032] = 16'h0000;
        rom[0][1033] = 16'h0000;
        rom[0][1034] = 16'h0000;
        rom[0][1035] = 16'h0000;
        rom[0][1036] = 16'h0000;
        rom[0][1037] = 16'h0000;
        rom[0][1038] = 16'h0000;
        rom[0][1039] = 16'h0000;
        rom[0][1040] = 16'h0000;
        rom[0][1041] = 16'h0000;
        rom[0][1042] = 16'h0000;
        rom[0][1043] = 16'h0000;
        rom[0][1044] = 16'h0000;
        rom[0][1045] = 16'h0000;
        rom[0][1046] = 16'h0000;
        rom[0][1047] = 16'h0000;
        rom[0][1048] = 16'h0000;
        rom[0][1049] = 16'h0000;
        rom[0][1050] = 16'h0000;
        rom[0][1051] = 16'h0000;
        rom[0][1052] = 16'h0000;
        rom[0][1053] = 16'h0000;
        rom[0][1054] = 16'h0000;
        rom[0][1055] = 16'h0000;
        rom[0][1056] = 16'h0000;
        rom[0][1057] = 16'h0000;
        rom[0][1058] = 16'h0000;
        rom[0][1059] = 16'h0000;
        rom[0][1060] = 16'h0000;
        rom[0][1061] = 16'h0000;
        rom[0][1062] = 16'h0000;
        rom[0][1063] = 16'h0000;
        rom[0][1064] = 16'h0000;
        rom[0][1065] = 16'h0000;
        rom[0][1066] = 16'h0000;
        rom[0][1067] = 16'h0000;
        rom[0][1068] = 16'h0000;
        rom[0][1069] = 16'h0000;
        rom[0][1070] = 16'h0000;
        rom[0][1071] = 16'h0000;
        rom[0][1072] = 16'h0000;
        rom[0][1073] = 16'h0000;
        rom[0][1074] = 16'h0000;
        rom[0][1075] = 16'h0000;
        rom[0][1076] = 16'h0000;
        rom[0][1077] = 16'h0000;
        rom[0][1078] = 16'h0065;
        rom[0][1079] = 16'hFFBF;
        rom[0][1080] = 16'hFFD5;
        rom[0][1081] = 16'hFFB8;
        rom[0][1082] = 16'hFFBF;
        rom[0][1083] = 16'hFF70;
        rom[0][1084] = 16'hFF12;
        rom[0][1085] = 16'hFF5A;
        rom[0][1086] = 16'hFFDC;
        rom[0][1087] = 16'hFFE3;
        rom[0][1088] = 16'hFFF9;
        rom[0][1089] = 16'hFFE3;
        rom[0][1090] = 16'h009F;
        rom[0][1091] = 16'h00AD;
        rom[0][1092] = 16'hFFE3;
        rom[0][1093] = 16'hFFDC;
        rom[0][1094] = 16'hFFCD;
        rom[0][1095] = 16'hFFA9;
        rom[0][1096] = 16'h000E;
        rom[0][1097] = 16'hFFA2;
        rom[0][1098] = 16'hFFF9;
        rom[0][1099] = 16'hFFC6;
        rom[0][1100] = 16'hFF77;
        rom[0][1101] = 16'hFEA6;
        rom[0][1102] = 16'hFE56;
        rom[0][1103] = 16'hFE73;
        rom[0][1104] = 16'hFF8D;
        rom[0][1105] = 16'hFF70;
        rom[0][1106] = 16'hFEC2;
        rom[0][1107] = 16'hFF20;
        rom[0][1108] = 16'hFF85;
        rom[0][1109] = 16'hFF20;
        rom[0][1110] = 16'h0000;
        rom[0][1111] = 16'h0000;
        rom[0][1112] = 16'h0000;
        rom[0][1113] = 16'h0000;
        rom[0][1114] = 16'h0000;
        rom[0][1115] = 16'h0000;
        rom[0][1116] = 16'h0000;
        rom[0][1117] = 16'h0000;
        rom[0][1118] = 16'h0000;
        rom[0][1119] = 16'h0000;
        rom[0][1120] = 16'h0000;
        rom[0][1121] = 16'h0000;
        rom[0][1122] = 16'h0000;
        rom[0][1123] = 16'h0000;
        rom[0][1124] = 16'h0000;
        rom[0][1125] = 16'h0000;
        rom[0][1126] = 16'h0000;
        rom[0][1127] = 16'h0000;
        rom[0][1128] = 16'h0000;
        rom[0][1129] = 16'h0000;
        rom[0][1130] = 16'h0000;
        rom[0][1131] = 16'h0000;
        rom[0][1132] = 16'h0000;
        rom[0][1133] = 16'h0000;
        rom[0][1134] = 16'h0000;
        rom[0][1135] = 16'h0000;
        rom[0][1136] = 16'h0000;
        rom[0][1137] = 16'h0000;
        rom[0][1138] = 16'h0000;
        rom[0][1139] = 16'h0000;
        rom[0][1140] = 16'h0000;
        rom[0][1141] = 16'h0000;
        rom[0][1142] = 16'h0000;
        rom[0][1143] = 16'h0000;
        rom[0][1144] = 16'h0000;
        rom[0][1145] = 16'h0000;
        rom[0][1146] = 16'h0000;
        rom[0][1147] = 16'h0000;
        rom[0][1148] = 16'h0000;
        rom[0][1149] = 16'h0000;
        rom[0][1150] = 16'h0000;
        rom[0][1151] = 16'h0000;
        rom[0][1152] = 16'h0000;
        rom[0][1153] = 16'h0000;
        rom[0][1154] = 16'h0000;
        rom[0][1155] = 16'h0000;
        rom[0][1156] = 16'h0000;
        rom[0][1157] = 16'h0000;
        rom[0][1158] = 16'h0000;
        rom[0][1159] = 16'h0000;
        rom[0][1160] = 16'h0000;
        rom[0][1161] = 16'h0000;
        rom[0][1162] = 16'h0000;
        rom[0][1163] = 16'h0000;
        rom[0][1164] = 16'h0000;
        rom[0][1165] = 16'h0000;
        rom[0][1166] = 16'h0000;
        rom[0][1167] = 16'h0000;
        rom[0][1168] = 16'h0000;
        rom[0][1169] = 16'h0000;
        rom[0][1170] = 16'h0000;
        rom[0][1171] = 16'h0000;
        rom[0][1172] = 16'h0000;
        rom[0][1173] = 16'h0000;
        rom[0][1174] = 16'h0000;
        rom[0][1175] = 16'h0000;
        rom[0][1176] = 16'h0194;
        rom[0][1177] = 16'h00F5;
        rom[0][1178] = 16'hFFC6;
        rom[0][1179] = 16'h0098;
        rom[0][1180] = 16'h0090;
        rom[0][1181] = 16'h004F;
        rom[0][1182] = 16'h00FD;
        rom[0][1183] = 16'h009F;
        rom[0][1184] = 16'h006C;
        rom[0][1185] = 16'h00AD;
        rom[0][1186] = 16'h00B4;
        rom[0][1187] = 16'h00AD;
        rom[0][1188] = 16'h00D9;
        rom[0][1189] = 16'h0089;
        rom[0][1190] = 16'h0057;
        rom[0][1191] = 16'h009F;
        rom[0][1192] = 16'h0041;
        rom[0][1193] = 16'h0016;
        rom[0][1194] = 16'h0007;
        rom[0][1195] = 16'hFEFC;
        rom[0][1196] = 16'hFF19;
        rom[0][1197] = 16'hFFB1;
        rom[0][1198] = 16'hFFDC;
        rom[0][1199] = 16'hFFA9;
        rom[0][1200] = 16'h0073;
        rom[0][1201] = 16'h00BC;
        rom[0][1202] = 16'h006C;
        rom[0][1203] = 16'h00D9;
        rom[0][1204] = 16'h00FD;
        rom[0][1205] = 16'h010B;
        rom[0][1206] = 16'h00C3;
        rom[0][1207] = 16'hFFC6;
        rom[0][1208] = 16'h0000;
        rom[0][1209] = 16'h0000;
        rom[0][1210] = 16'h0000;
        rom[0][1211] = 16'h0000;
        rom[0][1212] = 16'h0000;
        rom[0][1213] = 16'h0000;
        rom[0][1214] = 16'h0000;
        rom[0][1215] = 16'h0000;
        rom[0][1216] = 16'h0000;
        rom[0][1217] = 16'h0000;
        rom[0][1218] = 16'h0000;
        rom[0][1219] = 16'h0000;
        rom[0][1220] = 16'h0000;
        rom[0][1221] = 16'h0000;
        rom[0][1222] = 16'h0000;
        rom[0][1223] = 16'h0000;
        rom[0][1224] = 16'h0000;
        rom[0][1225] = 16'h0000;
        rom[0][1226] = 16'h0000;
        rom[0][1227] = 16'h0000;
        rom[0][1228] = 16'h0000;
        rom[0][1229] = 16'h0000;
        rom[0][1230] = 16'h0000;
        rom[0][1231] = 16'h0000;
        rom[0][1232] = 16'h0000;
        rom[0][1233] = 16'h0000;
        rom[0][1234] = 16'h0000;
        rom[0][1235] = 16'h0000;
        rom[0][1236] = 16'h0000;
        rom[0][1237] = 16'h0000;
        rom[0][1238] = 16'h0000;
        rom[0][1239] = 16'h0000;
        rom[0][1240] = 16'h0000;
        rom[0][1241] = 16'h0000;
        rom[0][1242] = 16'h0000;
        rom[0][1243] = 16'h0000;
        rom[0][1244] = 16'h0000;
        rom[0][1245] = 16'h0000;
        rom[0][1246] = 16'h0000;
        rom[0][1247] = 16'h0000;
        rom[0][1248] = 16'h0000;
        rom[0][1249] = 16'h0000;
        rom[0][1250] = 16'h0000;
        rom[0][1251] = 16'h0000;
        rom[0][1252] = 16'h0000;
        rom[0][1253] = 16'h0000;
        rom[0][1254] = 16'h0000;
        rom[0][1255] = 16'h0000;
        rom[0][1256] = 16'h0000;
        rom[0][1257] = 16'h0000;
        rom[0][1258] = 16'h0000;
        rom[0][1259] = 16'h0000;
        rom[0][1260] = 16'h0000;
        rom[0][1261] = 16'h0000;
        rom[0][1262] = 16'h0000;
        rom[0][1263] = 16'h0000;
        rom[0][1264] = 16'h0000;
        rom[0][1265] = 16'h0000;
        rom[0][1266] = 16'h0000;
        rom[0][1267] = 16'h0000;
        rom[0][1268] = 16'h0000;
        rom[0][1269] = 16'h0000;
        rom[0][1270] = 16'h0000;
        rom[0][1271] = 16'h0000;
        rom[0][1272] = 16'h0000;
        rom[0][1273] = 16'h0000;
        rom[1][0] = 16'h0082;
        rom[1][1] = 16'h0073;
        rom[1][2] = 16'h005E;
        rom[1][3] = 16'h003A;
        rom[1][4] = 16'h0016;
        rom[1][5] = 16'hFFF9;
        rom[1][6] = 16'h0119;
        rom[1][7] = 16'h017F;
        rom[1][8] = 16'h018D;
        rom[1][9] = 16'h017F;
        rom[1][10] = 16'h014C;
        rom[1][11] = 16'h00FD;
        rom[1][12] = 16'h00B4;
        rom[1][13] = 16'h0065;
        rom[1][14] = 16'hFFF9;
        rom[1][15] = 16'hFFA9;
        rom[1][16] = 16'hFF77;
        rom[1][17] = 16'hFF5A;
        rom[1][18] = 16'hFF44;
        rom[1][19] = 16'hFF3D;
        rom[1][20] = 16'hFF44;
        rom[1][21] = 16'hFF61;
        rom[1][22] = 16'hFF7E;
        rom[1][23] = 16'hFF94;
        rom[1][24] = 16'hFFB1;
        rom[1][25] = 16'hFFCD;
        rom[1][26] = 16'hFFEA;
        rom[1][27] = 16'h0007;
        rom[1][28] = 16'h002B;
        rom[1][29] = 16'h0041;
        rom[1][30] = 16'h005E;
        rom[1][31] = 16'h006C;
        rom[1][32] = 16'h0000;
        rom[1][33] = 16'h0000;
        rom[1][34] = 16'h0000;
        rom[1][35] = 16'h0000;
        rom[1][36] = 16'h0000;
        rom[1][37] = 16'h0000;
        rom[1][38] = 16'h0000;
        rom[1][39] = 16'h0000;
        rom[1][40] = 16'h0000;
        rom[1][41] = 16'h0000;
        rom[1][42] = 16'h0000;
        rom[1][43] = 16'h0000;
        rom[1][44] = 16'h0000;
        rom[1][45] = 16'h0000;
        rom[1][46] = 16'h0000;
        rom[1][47] = 16'h0000;
        rom[1][48] = 16'h0000;
        rom[1][49] = 16'h0000;
        rom[1][50] = 16'h0000;
        rom[1][51] = 16'h0000;
        rom[1][52] = 16'h0000;
        rom[1][53] = 16'h0000;
        rom[1][54] = 16'h0000;
        rom[1][55] = 16'h0000;
        rom[1][56] = 16'h0000;
        rom[1][57] = 16'h0000;
        rom[1][58] = 16'h0000;
        rom[1][59] = 16'h0000;
        rom[1][60] = 16'h0000;
        rom[1][61] = 16'h0000;
        rom[1][62] = 16'h0000;
        rom[1][63] = 16'h0000;
        rom[1][64] = 16'h0000;
        rom[1][65] = 16'h0000;
        rom[1][66] = 16'h0000;
        rom[1][67] = 16'h0000;
        rom[1][68] = 16'h0000;
        rom[1][69] = 16'h0000;
        rom[1][70] = 16'h0000;
        rom[1][71] = 16'h0000;
        rom[1][72] = 16'h0000;
        rom[1][73] = 16'h0000;
        rom[1][74] = 16'h0000;
        rom[1][75] = 16'h0000;
        rom[1][76] = 16'h0000;
        rom[1][77] = 16'h0000;
        rom[1][78] = 16'h0000;
        rom[1][79] = 16'h0000;
        rom[1][80] = 16'h0000;
        rom[1][81] = 16'h0000;
        rom[1][82] = 16'h0000;
        rom[1][83] = 16'h0000;
        rom[1][84] = 16'h0000;
        rom[1][85] = 16'h0000;
        rom[1][86] = 16'h0000;
        rom[1][87] = 16'h0000;
        rom[1][88] = 16'h0000;
        rom[1][89] = 16'h0000;
        rom[1][90] = 16'h0000;
        rom[1][91] = 16'h0000;
        rom[1][92] = 16'h0000;
        rom[1][93] = 16'h0000;
        rom[1][94] = 16'h0000;
        rom[1][95] = 16'h0000;
        rom[1][96] = 16'h0000;
        rom[1][97] = 16'h0000;
        rom[1][98] = 16'h00FD;
        rom[1][99] = 16'h00C3;
        rom[1][100] = 16'h00AD;
        rom[1][101] = 16'h007B;
        rom[1][102] = 16'h004F;
        rom[1][103] = 16'h003A;
        rom[1][104] = 16'h009F;
        rom[1][105] = 16'h00BC;
        rom[1][106] = 16'h00AD;
        rom[1][107] = 16'h0098;
        rom[1][108] = 16'h007B;
        rom[1][109] = 16'h005E;
        rom[1][110] = 16'h0065;
        rom[1][111] = 16'h006C;
        rom[1][112] = 16'h0073;
        rom[1][113] = 16'h0090;
        rom[1][114] = 16'h007B;
        rom[1][115] = 16'h0048;
        rom[1][116] = 16'h000E;
        rom[1][117] = 16'hFFE3;
        rom[1][118] = 16'hFFBF;
        rom[1][119] = 16'hFFC6;
        rom[1][120] = 16'hFFDC;
        rom[1][121] = 16'hFFF2;
        rom[1][122] = 16'h0007;
        rom[1][123] = 16'h0007;
        rom[1][124] = 16'h0016;
        rom[1][125] = 16'h0033;
        rom[1][126] = 16'h004F;
        rom[1][127] = 16'h0065;
        rom[1][128] = 16'h007B;
        rom[1][129] = 16'h00AD;
        rom[1][130] = 16'h0000;
        rom[1][131] = 16'h0000;
        rom[1][132] = 16'h0000;
        rom[1][133] = 16'h0000;
        rom[1][134] = 16'h0000;
        rom[1][135] = 16'h0000;
        rom[1][136] = 16'h0000;
        rom[1][137] = 16'h0000;
        rom[1][138] = 16'h0000;
        rom[1][139] = 16'h0000;
        rom[1][140] = 16'h0000;
        rom[1][141] = 16'h0000;
        rom[1][142] = 16'h0000;
        rom[1][143] = 16'h0000;
        rom[1][144] = 16'h0000;
        rom[1][145] = 16'h0000;
        rom[1][146] = 16'h0000;
        rom[1][147] = 16'h0000;
        rom[1][148] = 16'h0000;
        rom[1][149] = 16'h0000;
        rom[1][150] = 16'h0000;
        rom[1][151] = 16'h0000;
        rom[1][152] = 16'h0000;
        rom[1][153] = 16'h0000;
        rom[1][154] = 16'h0000;
        rom[1][155] = 16'h0000;
        rom[1][156] = 16'h0000;
        rom[1][157] = 16'h0000;
        rom[1][158] = 16'h0000;
        rom[1][159] = 16'h0000;
        rom[1][160] = 16'h0000;
        rom[1][161] = 16'h0000;
        rom[1][162] = 16'h0000;
        rom[1][163] = 16'h0000;
        rom[1][164] = 16'h0000;
        rom[1][165] = 16'h0000;
        rom[1][166] = 16'h0000;
        rom[1][167] = 16'h0000;
        rom[1][168] = 16'h0000;
        rom[1][169] = 16'h0000;
        rom[1][170] = 16'h0000;
        rom[1][171] = 16'h0000;
        rom[1][172] = 16'h0000;
        rom[1][173] = 16'h0000;
        rom[1][174] = 16'h0000;
        rom[1][175] = 16'h0000;
        rom[1][176] = 16'h0000;
        rom[1][177] = 16'h0000;
        rom[1][178] = 16'h0000;
        rom[1][179] = 16'h0000;
        rom[1][180] = 16'h0000;
        rom[1][181] = 16'h0000;
        rom[1][182] = 16'h0000;
        rom[1][183] = 16'h0000;
        rom[1][184] = 16'h0000;
        rom[1][185] = 16'h0000;
        rom[1][186] = 16'h0000;
        rom[1][187] = 16'h0000;
        rom[1][188] = 16'h0000;
        rom[1][189] = 16'h0000;
        rom[1][190] = 16'h0000;
        rom[1][191] = 16'h0000;
        rom[1][192] = 16'h0000;
        rom[1][193] = 16'h0000;
        rom[1][194] = 16'h0000;
        rom[1][195] = 16'h0000;
        rom[1][196] = 16'h0065;
        rom[1][197] = 16'h0048;
        rom[1][198] = 16'h0041;
        rom[1][199] = 16'h002B;
        rom[1][200] = 16'h003A;
        rom[1][201] = 16'h001D;
        rom[1][202] = 16'hFECA;
        rom[1][203] = 16'hFF36;
        rom[1][204] = 16'hFF20;
        rom[1][205] = 16'hFED8;
        rom[1][206] = 16'hFEEE;
        rom[1][207] = 16'hFF61;
        rom[1][208] = 16'hFFC6;
        rom[1][209] = 16'h000E;
        rom[1][210] = 16'h009F;
        rom[1][211] = 16'h00FD;
        rom[1][212] = 16'h0112;
        rom[1][213] = 16'h00D1;
        rom[1][214] = 16'h009F;
        rom[1][215] = 16'h007B;
        rom[1][216] = 16'h006C;
        rom[1][217] = 16'h005E;
        rom[1][218] = 16'h005E;
        rom[1][219] = 16'h007B;
        rom[1][220] = 16'h0073;
        rom[1][221] = 16'h004F;
        rom[1][222] = 16'h0041;
        rom[1][223] = 16'h002B;
        rom[1][224] = 16'h002B;
        rom[1][225] = 16'h0065;
        rom[1][226] = 16'h006C;
        rom[1][227] = 16'h0073;
        rom[1][228] = 16'h0000;
        rom[1][229] = 16'h0000;
        rom[1][230] = 16'h0000;
        rom[1][231] = 16'h0000;
        rom[1][232] = 16'h0000;
        rom[1][233] = 16'h0000;
        rom[1][234] = 16'h0000;
        rom[1][235] = 16'h0000;
        rom[1][236] = 16'h0000;
        rom[1][237] = 16'h0000;
        rom[1][238] = 16'h0000;
        rom[1][239] = 16'h0000;
        rom[1][240] = 16'h0000;
        rom[1][241] = 16'h0000;
        rom[1][242] = 16'h0000;
        rom[1][243] = 16'h0000;
        rom[1][244] = 16'h0000;
        rom[1][245] = 16'h0000;
        rom[1][246] = 16'h0000;
        rom[1][247] = 16'h0000;
        rom[1][248] = 16'h0000;
        rom[1][249] = 16'h0000;
        rom[1][250] = 16'h0000;
        rom[1][251] = 16'h0000;
        rom[1][252] = 16'h0000;
        rom[1][253] = 16'h0000;
        rom[1][254] = 16'h0000;
        rom[1][255] = 16'h0000;
        rom[1][256] = 16'h0000;
        rom[1][257] = 16'h0000;
        rom[1][258] = 16'h0000;
        rom[1][259] = 16'h0000;
        rom[1][260] = 16'h0000;
        rom[1][261] = 16'h0000;
        rom[1][262] = 16'h0000;
        rom[1][263] = 16'h0000;
        rom[1][264] = 16'h0000;
        rom[1][265] = 16'h0000;
        rom[1][266] = 16'h0000;
        rom[1][267] = 16'h0000;
        rom[1][268] = 16'h0000;
        rom[1][269] = 16'h0000;
        rom[1][270] = 16'h0000;
        rom[1][271] = 16'h0000;
        rom[1][272] = 16'h0000;
        rom[1][273] = 16'h0000;
        rom[1][274] = 16'h0000;
        rom[1][275] = 16'h0000;
        rom[1][276] = 16'h0000;
        rom[1][277] = 16'h0000;
        rom[1][278] = 16'h0000;
        rom[1][279] = 16'h0000;
        rom[1][280] = 16'h0000;
        rom[1][281] = 16'h0000;
        rom[1][282] = 16'h0000;
        rom[1][283] = 16'h0000;
        rom[1][284] = 16'h0000;
        rom[1][285] = 16'h0000;
        rom[1][286] = 16'h0000;
        rom[1][287] = 16'h0000;
        rom[1][288] = 16'h0000;
        rom[1][289] = 16'h0000;
        rom[1][290] = 16'h0000;
        rom[1][291] = 16'h0000;
        rom[1][292] = 16'h0000;
        rom[1][293] = 16'h0000;
        rom[1][294] = 16'h00D9;
        rom[1][295] = 16'h00D1;
        rom[1][296] = 16'h00BC;
        rom[1][297] = 16'h009F;
        rom[1][298] = 16'h009F;
        rom[1][299] = 16'h0048;
        rom[1][300] = 16'hFF4C;
        rom[1][301] = 16'hFFB1;
        rom[1][302] = 16'h002B;
        rom[1][303] = 16'hFFEA;
        rom[1][304] = 16'hFF8D;
        rom[1][305] = 16'hFF77;
        rom[1][306] = 16'hFF77;
        rom[1][307] = 16'hFF77;
        rom[1][308] = 16'hFFB1;
        rom[1][309] = 16'h000E;
        rom[1][310] = 16'h0041;
        rom[1][311] = 16'h0033;
        rom[1][312] = 16'h0057;
        rom[1][313] = 16'h0057;
        rom[1][314] = 16'h007B;
        rom[1][315] = 16'h0098;
        rom[1][316] = 16'h009F;
        rom[1][317] = 16'h00BC;
        rom[1][318] = 16'h00E0;
        rom[1][319] = 16'h00CA;
        rom[1][320] = 16'h00CA;
        rom[1][321] = 16'h00D1;
        rom[1][322] = 16'h00E0;
        rom[1][323] = 16'h0119;
        rom[1][324] = 16'h0119;
        rom[1][325] = 16'h0104;
        rom[1][326] = 16'h0000;
        rom[1][327] = 16'h0000;
        rom[1][328] = 16'h0000;
        rom[1][329] = 16'h0000;
        rom[1][330] = 16'h0000;
        rom[1][331] = 16'h0000;
        rom[1][332] = 16'h0000;
        rom[1][333] = 16'h0000;
        rom[1][334] = 16'h0000;
        rom[1][335] = 16'h0000;
        rom[1][336] = 16'h0000;
        rom[1][337] = 16'h0000;
        rom[1][338] = 16'h0000;
        rom[1][339] = 16'h0000;
        rom[1][340] = 16'h0000;
        rom[1][341] = 16'h0000;
        rom[1][342] = 16'h0000;
        rom[1][343] = 16'h0000;
        rom[1][344] = 16'h0000;
        rom[1][345] = 16'h0000;
        rom[1][346] = 16'h0000;
        rom[1][347] = 16'h0000;
        rom[1][348] = 16'h0000;
        rom[1][349] = 16'h0000;
        rom[1][350] = 16'h0000;
        rom[1][351] = 16'h0000;
        rom[1][352] = 16'h0000;
        rom[1][353] = 16'h0000;
        rom[1][354] = 16'h0000;
        rom[1][355] = 16'h0000;
        rom[1][356] = 16'h0000;
        rom[1][357] = 16'h0000;
        rom[1][358] = 16'h0000;
        rom[1][359] = 16'h0000;
        rom[1][360] = 16'h0000;
        rom[1][361] = 16'h0000;
        rom[1][362] = 16'h0000;
        rom[1][363] = 16'h0000;
        rom[1][364] = 16'h0000;
        rom[1][365] = 16'h0000;
        rom[1][366] = 16'h0000;
        rom[1][367] = 16'h0000;
        rom[1][368] = 16'h0000;
        rom[1][369] = 16'h0000;
        rom[1][370] = 16'h0000;
        rom[1][371] = 16'h0000;
        rom[1][372] = 16'h0000;
        rom[1][373] = 16'h0000;
        rom[1][374] = 16'h0000;
        rom[1][375] = 16'h0000;
        rom[1][376] = 16'h0000;
        rom[1][377] = 16'h0000;
        rom[1][378] = 16'h0000;
        rom[1][379] = 16'h0000;
        rom[1][380] = 16'h0000;
        rom[1][381] = 16'h0000;
        rom[1][382] = 16'h0000;
        rom[1][383] = 16'h0000;
        rom[1][384] = 16'h0000;
        rom[1][385] = 16'h0000;
        rom[1][386] = 16'h0000;
        rom[1][387] = 16'h0000;
        rom[1][388] = 16'h0000;
        rom[1][389] = 16'h0000;
        rom[1][390] = 16'h0000;
        rom[1][391] = 16'h0000;
        rom[1][392] = 16'h0007;
        rom[1][393] = 16'h0057;
        rom[1][394] = 16'h007B;
        rom[1][395] = 16'h0098;
        rom[1][396] = 16'h0073;
        rom[1][397] = 16'h004F;
        rom[1][398] = 16'hFFE3;
        rom[1][399] = 16'hFF7E;
        rom[1][400] = 16'hFEAD;
        rom[1][401] = 16'hFE5D;
        rom[1][402] = 16'hFE7A;
        rom[1][403] = 16'hFEA6;
        rom[1][404] = 16'hFECA;
        rom[1][405] = 16'hFED8;
        rom[1][406] = 16'hFEFC;
        rom[1][407] = 16'hFF4C;
        rom[1][408] = 16'hFFD5;
        rom[1][409] = 16'h004F;
        rom[1][410] = 16'h00CA;
        rom[1][411] = 16'h00C3;
        rom[1][412] = 16'h009F;
        rom[1][413] = 16'h00C3;
        rom[1][414] = 16'h00D1;
        rom[1][415] = 16'h00C3;
        rom[1][416] = 16'h00CA;
        rom[1][417] = 16'h00D9;
        rom[1][418] = 16'h0098;
        rom[1][419] = 16'h007B;
        rom[1][420] = 16'h0073;
        rom[1][421] = 16'h0073;
        rom[1][422] = 16'h004F;
        rom[1][423] = 16'h0057;
        rom[1][424] = 16'h0000;
        rom[1][425] = 16'h0000;
        rom[1][426] = 16'h0000;
        rom[1][427] = 16'h0000;
        rom[1][428] = 16'h0000;
        rom[1][429] = 16'h0000;
        rom[1][430] = 16'h0000;
        rom[1][431] = 16'h0000;
        rom[1][432] = 16'h0000;
        rom[1][433] = 16'h0000;
        rom[1][434] = 16'h0000;
        rom[1][435] = 16'h0000;
        rom[1][436] = 16'h0000;
        rom[1][437] = 16'h0000;
        rom[1][438] = 16'h0000;
        rom[1][439] = 16'h0000;
        rom[1][440] = 16'h0000;
        rom[1][441] = 16'h0000;
        rom[1][442] = 16'h0000;
        rom[1][443] = 16'h0000;
        rom[1][444] = 16'h0000;
        rom[1][445] = 16'h0000;
        rom[1][446] = 16'h0000;
        rom[1][447] = 16'h0000;
        rom[1][448] = 16'h0000;
        rom[1][449] = 16'h0000;
        rom[1][450] = 16'h0000;
        rom[1][451] = 16'h0000;
        rom[1][452] = 16'h0000;
        rom[1][453] = 16'h0000;
        rom[1][454] = 16'h0000;
        rom[1][455] = 16'h0000;
        rom[1][456] = 16'h0000;
        rom[1][457] = 16'h0000;
        rom[1][458] = 16'h0000;
        rom[1][459] = 16'h0000;
        rom[1][460] = 16'h0000;
        rom[1][461] = 16'h0000;
        rom[1][462] = 16'h0000;
        rom[1][463] = 16'h0000;
        rom[1][464] = 16'h0000;
        rom[1][465] = 16'h0000;
        rom[1][466] = 16'h0000;
        rom[1][467] = 16'h0000;
        rom[1][468] = 16'h0000;
        rom[1][469] = 16'h0000;
        rom[1][470] = 16'h0000;
        rom[1][471] = 16'h0000;
        rom[1][472] = 16'h0000;
        rom[1][473] = 16'h0000;
        rom[1][474] = 16'h0000;
        rom[1][475] = 16'h0000;
        rom[1][476] = 16'h0000;
        rom[1][477] = 16'h0000;
        rom[1][478] = 16'h0000;
        rom[1][479] = 16'h0000;
        rom[1][480] = 16'h0000;
        rom[1][481] = 16'h0000;
        rom[1][482] = 16'h0000;
        rom[1][483] = 16'h0000;
        rom[1][484] = 16'h0000;
        rom[1][485] = 16'h0000;
        rom[1][486] = 16'h0000;
        rom[1][487] = 16'h0000;
        rom[1][488] = 16'h0000;
        rom[1][489] = 16'h0000;
        rom[1][490] = 16'h00BC;
        rom[1][491] = 16'h00E7;
        rom[1][492] = 16'h00D1;
        rom[1][493] = 16'h00CA;
        rom[1][494] = 16'h00AD;
        rom[1][495] = 16'h00E0;
        rom[1][496] = 16'h0208;
        rom[1][497] = 16'h01D5;
        rom[1][498] = 16'h014C;
        rom[1][499] = 16'h0119;
        rom[1][500] = 16'h0162;
        rom[1][501] = 16'h01DC;
        rom[1][502] = 16'h01F9;
        rom[1][503] = 16'h0200;
        rom[1][504] = 16'h01D5;
        rom[1][505] = 16'h00D1;
        rom[1][506] = 16'h0048;
        rom[1][507] = 16'h00BC;
        rom[1][508] = 16'h00FD;
        rom[1][509] = 16'h00F5;
        rom[1][510] = 16'h00A6;
        rom[1][511] = 16'h00C3;
        rom[1][512] = 16'h00FD;
        rom[1][513] = 16'h0104;
        rom[1][514] = 16'h00F5;
        rom[1][515] = 16'h010B;
        rom[1][516] = 16'h00E7;
        rom[1][517] = 16'h00AD;
        rom[1][518] = 16'h0089;
        rom[1][519] = 16'h00C3;
        rom[1][520] = 16'h010B;
        rom[1][521] = 16'h010B;
        rom[1][522] = 16'h0000;
        rom[1][523] = 16'h0000;
        rom[1][524] = 16'h0000;
        rom[1][525] = 16'h0000;
        rom[1][526] = 16'h0000;
        rom[1][527] = 16'h0000;
        rom[1][528] = 16'h0000;
        rom[1][529] = 16'h0000;
        rom[1][530] = 16'h0000;
        rom[1][531] = 16'h0000;
        rom[1][532] = 16'h0000;
        rom[1][533] = 16'h0000;
        rom[1][534] = 16'h0000;
        rom[1][535] = 16'h0000;
        rom[1][536] = 16'h0000;
        rom[1][537] = 16'h0000;
        rom[1][538] = 16'h0000;
        rom[1][539] = 16'h0000;
        rom[1][540] = 16'h0000;
        rom[1][541] = 16'h0000;
        rom[1][542] = 16'h0000;
        rom[1][543] = 16'h0000;
        rom[1][544] = 16'h0000;
        rom[1][545] = 16'h0000;
        rom[1][546] = 16'h0000;
        rom[1][547] = 16'h0000;
        rom[1][548] = 16'h0000;
        rom[1][549] = 16'h0000;
        rom[1][550] = 16'h0000;
        rom[1][551] = 16'h0000;
        rom[1][552] = 16'h0000;
        rom[1][553] = 16'h0000;
        rom[1][554] = 16'h0000;
        rom[1][555] = 16'h0000;
        rom[1][556] = 16'h0000;
        rom[1][557] = 16'h0000;
        rom[1][558] = 16'h0000;
        rom[1][559] = 16'h0000;
        rom[1][560] = 16'h0000;
        rom[1][561] = 16'h0000;
        rom[1][562] = 16'h0000;
        rom[1][563] = 16'h0000;
        rom[1][564] = 16'h0000;
        rom[1][565] = 16'h0000;
        rom[1][566] = 16'h0000;
        rom[1][567] = 16'h0000;
        rom[1][568] = 16'h0000;
        rom[1][569] = 16'h0000;
        rom[1][570] = 16'h0000;
        rom[1][571] = 16'h0000;
        rom[1][572] = 16'h0000;
        rom[1][573] = 16'h0000;
        rom[1][574] = 16'h0000;
        rom[1][575] = 16'h0000;
        rom[1][576] = 16'h0000;
        rom[1][577] = 16'h0000;
        rom[1][578] = 16'h0000;
        rom[1][579] = 16'h0000;
        rom[1][580] = 16'h0000;
        rom[1][581] = 16'h0000;
        rom[1][582] = 16'h0000;
        rom[1][583] = 16'h0000;
        rom[1][584] = 16'h0000;
        rom[1][585] = 16'h0000;
        rom[1][586] = 16'h0000;
        rom[1][587] = 16'h0000;
        rom[1][588] = 16'h00C3;
        rom[1][589] = 16'h009F;
        rom[1][590] = 16'h0065;
        rom[1][591] = 16'h004F;
        rom[1][592] = 16'h0082;
        rom[1][593] = 16'h00BC;
        rom[1][594] = 16'hFE90;
        rom[1][595] = 16'hFE1C;
        rom[1][596] = 16'hFE1C;
        rom[1][597] = 16'hFE7A;
        rom[1][598] = 16'hFED1;
        rom[1][599] = 16'hFF2F;
        rom[1][600] = 16'hFF94;
        rom[1][601] = 16'h001D;
        rom[1][602] = 16'h0098;
        rom[1][603] = 16'h0082;
        rom[1][604] = 16'h0048;
        rom[1][605] = 16'h0089;
        rom[1][606] = 16'h00D9;
        rom[1][607] = 16'h0104;
        rom[1][608] = 16'h00B4;
        rom[1][609] = 16'h007B;
        rom[1][610] = 16'h0090;
        rom[1][611] = 16'h009F;
        rom[1][612] = 16'h00A6;
        rom[1][613] = 16'h00C3;
        rom[1][614] = 16'h00E7;
        rom[1][615] = 16'h00D1;
        rom[1][616] = 16'h006C;
        rom[1][617] = 16'h0098;
        rom[1][618] = 16'h00FD;
        rom[1][619] = 16'h00F5;
        rom[1][620] = 16'h0000;
        rom[1][621] = 16'h0000;
        rom[1][622] = 16'h0000;
        rom[1][623] = 16'h0000;
        rom[1][624] = 16'h0000;
        rom[1][625] = 16'h0000;
        rom[1][626] = 16'h0000;
        rom[1][627] = 16'h0000;
        rom[1][628] = 16'h0000;
        rom[1][629] = 16'h0000;
        rom[1][630] = 16'h0000;
        rom[1][631] = 16'h0000;
        rom[1][632] = 16'h0000;
        rom[1][633] = 16'h0000;
        rom[1][634] = 16'h0000;
        rom[1][635] = 16'h0000;
        rom[1][636] = 16'h0000;
        rom[1][637] = 16'h0000;
        rom[1][638] = 16'h0000;
        rom[1][639] = 16'h0000;
        rom[1][640] = 16'h0000;
        rom[1][641] = 16'h0000;
        rom[1][642] = 16'h0000;
        rom[1][643] = 16'h0000;
        rom[1][644] = 16'h0000;
        rom[1][645] = 16'h0000;
        rom[1][646] = 16'h0000;
        rom[1][647] = 16'h0000;
        rom[1][648] = 16'h0000;
        rom[1][649] = 16'h0000;
        rom[1][650] = 16'h0000;
        rom[1][651] = 16'h0000;
        rom[1][652] = 16'h0000;
        rom[1][653] = 16'h0000;
        rom[1][654] = 16'h0000;
        rom[1][655] = 16'h0000;
        rom[1][656] = 16'h0000;
        rom[1][657] = 16'h0000;
        rom[1][658] = 16'h0000;
        rom[1][659] = 16'h0000;
        rom[1][660] = 16'h0000;
        rom[1][661] = 16'h0000;
        rom[1][662] = 16'h0000;
        rom[1][663] = 16'h0000;
        rom[1][664] = 16'h0000;
        rom[1][665] = 16'h0000;
        rom[1][666] = 16'h0000;
        rom[1][667] = 16'h0000;
        rom[1][668] = 16'h0000;
        rom[1][669] = 16'h0000;
        rom[1][670] = 16'h0000;
        rom[1][671] = 16'h0000;
        rom[1][672] = 16'h0000;
        rom[1][673] = 16'h0000;
        rom[1][674] = 16'h0000;
        rom[1][675] = 16'h0000;
        rom[1][676] = 16'h0000;
        rom[1][677] = 16'h0000;
        rom[1][678] = 16'h0000;
        rom[1][679] = 16'h0000;
        rom[1][680] = 16'h0000;
        rom[1][681] = 16'h0000;
        rom[1][682] = 16'h0000;
        rom[1][683] = 16'h0000;
        rom[1][684] = 16'h0000;
        rom[1][685] = 16'h0000;
        rom[1][686] = 16'h00AD;
        rom[1][687] = 16'h00D1;
        rom[1][688] = 16'h0121;
        rom[1][689] = 16'h0112;
        rom[1][690] = 16'h0119;
        rom[1][691] = 16'h00F5;
        rom[1][692] = 16'h003A;
        rom[1][693] = 16'hFFE3;
        rom[1][694] = 16'h001D;
        rom[1][695] = 16'h0089;
        rom[1][696] = 16'h00CA;
        rom[1][697] = 16'h00E0;
        rom[1][698] = 16'h00A6;
        rom[1][699] = 16'h009F;
        rom[1][700] = 16'h010B;
        rom[1][701] = 16'h015A;
        rom[1][702] = 16'h0145;
        rom[1][703] = 16'h00E7;
        rom[1][704] = 16'h00C3;
        rom[1][705] = 16'h0104;
        rom[1][706] = 16'h010B;
        rom[1][707] = 16'h00F5;
        rom[1][708] = 16'h00E0;
        rom[1][709] = 16'h00D9;
        rom[1][710] = 16'h00CA;
        rom[1][711] = 16'h0119;
        rom[1][712] = 16'h0136;
        rom[1][713] = 16'h010B;
        rom[1][714] = 16'h0112;
        rom[1][715] = 16'h00FD;
        rom[1][716] = 16'h010B;
        rom[1][717] = 16'h00E0;
        rom[1][718] = 16'h0000;
        rom[1][719] = 16'h0000;
        rom[1][720] = 16'h0000;
        rom[1][721] = 16'h0000;
        rom[1][722] = 16'h0000;
        rom[1][723] = 16'h0000;
        rom[1][724] = 16'h0000;
        rom[1][725] = 16'h0000;
        rom[1][726] = 16'h0000;
        rom[1][727] = 16'h0000;
        rom[1][728] = 16'h0000;
        rom[1][729] = 16'h0000;
        rom[1][730] = 16'h0000;
        rom[1][731] = 16'h0000;
        rom[1][732] = 16'h0000;
        rom[1][733] = 16'h0000;
        rom[1][734] = 16'h0000;
        rom[1][735] = 16'h0000;
        rom[1][736] = 16'h0000;
        rom[1][737] = 16'h0000;
        rom[1][738] = 16'h0000;
        rom[1][739] = 16'h0000;
        rom[1][740] = 16'h0000;
        rom[1][741] = 16'h0000;
        rom[1][742] = 16'h0000;
        rom[1][743] = 16'h0000;
        rom[1][744] = 16'h0000;
        rom[1][745] = 16'h0000;
        rom[1][746] = 16'h0000;
        rom[1][747] = 16'h0000;
        rom[1][748] = 16'h0000;
        rom[1][749] = 16'h0000;
        rom[1][750] = 16'h0000;
        rom[1][751] = 16'h0000;
        rom[1][752] = 16'h0000;
        rom[1][753] = 16'h0000;
        rom[1][754] = 16'h0000;
        rom[1][755] = 16'h0000;
        rom[1][756] = 16'h0000;
        rom[1][757] = 16'h0000;
        rom[1][758] = 16'h0000;
        rom[1][759] = 16'h0000;
        rom[1][760] = 16'h0000;
        rom[1][761] = 16'h0000;
        rom[1][762] = 16'h0000;
        rom[1][763] = 16'h0000;
        rom[1][764] = 16'h0000;
        rom[1][765] = 16'h0000;
        rom[1][766] = 16'h0000;
        rom[1][767] = 16'h0000;
        rom[1][768] = 16'h0000;
        rom[1][769] = 16'h0000;
        rom[1][770] = 16'h0000;
        rom[1][771] = 16'h0000;
        rom[1][772] = 16'h0000;
        rom[1][773] = 16'h0000;
        rom[1][774] = 16'h0000;
        rom[1][775] = 16'h0000;
        rom[1][776] = 16'h0000;
        rom[1][777] = 16'h0000;
        rom[1][778] = 16'h0000;
        rom[1][779] = 16'h0000;
        rom[1][780] = 16'h0000;
        rom[1][781] = 16'h0000;
        rom[1][782] = 16'h0000;
        rom[1][783] = 16'h0000;
        rom[1][784] = 16'h0098;
        rom[1][785] = 16'h00EE;
        rom[1][786] = 16'h00E7;
        rom[1][787] = 16'h0104;
        rom[1][788] = 16'h00BC;
        rom[1][789] = 16'h0082;
        rom[1][790] = 16'hFF61;
        rom[1][791] = 16'hFF3D;
        rom[1][792] = 16'hFFB1;
        rom[1][793] = 16'h0000;
        rom[1][794] = 16'h000E;
        rom[1][795] = 16'hFFB8;
        rom[1][796] = 16'hFF85;
        rom[1][797] = 16'hFF53;
        rom[1][798] = 16'hFFA2;
        rom[1][799] = 16'h0057;
        rom[1][800] = 16'h00F5;
        rom[1][801] = 16'h00B4;
        rom[1][802] = 16'h003A;
        rom[1][803] = 16'h00B4;
        rom[1][804] = 16'h0098;
        rom[1][805] = 16'h0089;
        rom[1][806] = 16'h00A6;
        rom[1][807] = 16'h0089;
        rom[1][808] = 16'h0090;
        rom[1][809] = 16'h00E7;
        rom[1][810] = 16'h0104;
        rom[1][811] = 16'h0082;
        rom[1][812] = 16'h009F;
        rom[1][813] = 16'h0090;
        rom[1][814] = 16'h0089;
        rom[1][815] = 16'h0033;
        rom[1][816] = 16'h0000;
        rom[1][817] = 16'h0000;
        rom[1][818] = 16'h0000;
        rom[1][819] = 16'h0000;
        rom[1][820] = 16'h0000;
        rom[1][821] = 16'h0000;
        rom[1][822] = 16'h0000;
        rom[1][823] = 16'h0000;
        rom[1][824] = 16'h0000;
        rom[1][825] = 16'h0000;
        rom[1][826] = 16'h0000;
        rom[1][827] = 16'h0000;
        rom[1][828] = 16'h0000;
        rom[1][829] = 16'h0000;
        rom[1][830] = 16'h0000;
        rom[1][831] = 16'h0000;
        rom[1][832] = 16'h0000;
        rom[1][833] = 16'h0000;
        rom[1][834] = 16'h0000;
        rom[1][835] = 16'h0000;
        rom[1][836] = 16'h0000;
        rom[1][837] = 16'h0000;
        rom[1][838] = 16'h0000;
        rom[1][839] = 16'h0000;
        rom[1][840] = 16'h0000;
        rom[1][841] = 16'h0000;
        rom[1][842] = 16'h0000;
        rom[1][843] = 16'h0000;
        rom[1][844] = 16'h0000;
        rom[1][845] = 16'h0000;
        rom[1][846] = 16'h0000;
        rom[1][847] = 16'h0000;
        rom[1][848] = 16'h0000;
        rom[1][849] = 16'h0000;
        rom[1][850] = 16'h0000;
        rom[1][851] = 16'h0000;
        rom[1][852] = 16'h0000;
        rom[1][853] = 16'h0000;
        rom[1][854] = 16'h0000;
        rom[1][855] = 16'h0000;
        rom[1][856] = 16'h0000;
        rom[1][857] = 16'h0000;
        rom[1][858] = 16'h0000;
        rom[1][859] = 16'h0000;
        rom[1][860] = 16'h0000;
        rom[1][861] = 16'h0000;
        rom[1][862] = 16'h0000;
        rom[1][863] = 16'h0000;
        rom[1][864] = 16'h0000;
        rom[1][865] = 16'h0000;
        rom[1][866] = 16'h0000;
        rom[1][867] = 16'h0000;
        rom[1][868] = 16'h0000;
        rom[1][869] = 16'h0000;
        rom[1][870] = 16'h0000;
        rom[1][871] = 16'h0000;
        rom[1][872] = 16'h0000;
        rom[1][873] = 16'h0000;
        rom[1][874] = 16'h0000;
        rom[1][875] = 16'h0000;
        rom[1][876] = 16'h0000;
        rom[1][877] = 16'h0000;
        rom[1][878] = 16'h0000;
        rom[1][879] = 16'h0000;
        rom[1][880] = 16'h0000;
        rom[1][881] = 16'h0000;
        rom[1][882] = 16'h01B8;
        rom[1][883] = 16'h01B1;
        rom[1][884] = 16'h00EE;
        rom[1][885] = 16'h00FD;
        rom[1][886] = 16'h00E0;
        rom[1][887] = 16'h0136;
        rom[1][888] = 16'h02A6;
        rom[1][889] = 16'h0225;
        rom[1][890] = 16'h0194;
        rom[1][891] = 16'h019B;
        rom[1][892] = 16'h01DC;
        rom[1][893] = 16'h01EB;
        rom[1][894] = 16'h01EB;
        rom[1][895] = 16'h0128;
        rom[1][896] = 16'h0007;
        rom[1][897] = 16'hFFB1;
        rom[1][898] = 16'h001D;
        rom[1][899] = 16'h0048;
        rom[1][900] = 16'h0098;
        rom[1][901] = 16'h0112;
        rom[1][902] = 16'h00B4;
        rom[1][903] = 16'h0073;
        rom[1][904] = 16'h00C3;
        rom[1][905] = 16'h00EE;
        rom[1][906] = 16'h0119;
        rom[1][907] = 16'h0128;
        rom[1][908] = 16'h00D1;
        rom[1][909] = 16'h00AD;
        rom[1][910] = 16'h00E7;
        rom[1][911] = 16'h010B;
        rom[1][912] = 16'h0136;
        rom[1][913] = 16'h0121;
        rom[1][914] = 16'h0000;
        rom[1][915] = 16'h0000;
        rom[1][916] = 16'h0000;
        rom[1][917] = 16'h0000;
        rom[1][918] = 16'h0000;
        rom[1][919] = 16'h0000;
        rom[1][920] = 16'h0000;
        rom[1][921] = 16'h0000;
        rom[1][922] = 16'h0000;
        rom[1][923] = 16'h0000;
        rom[1][924] = 16'h0000;
        rom[1][925] = 16'h0000;
        rom[1][926] = 16'h0000;
        rom[1][927] = 16'h0000;
        rom[1][928] = 16'h0000;
        rom[1][929] = 16'h0000;
        rom[1][930] = 16'h0000;
        rom[1][931] = 16'h0000;
        rom[1][932] = 16'h0000;
        rom[1][933] = 16'h0000;
        rom[1][934] = 16'h0000;
        rom[1][935] = 16'h0000;
        rom[1][936] = 16'h0000;
        rom[1][937] = 16'h0000;
        rom[1][938] = 16'h0000;
        rom[1][939] = 16'h0000;
        rom[1][940] = 16'h0000;
        rom[1][941] = 16'h0000;
        rom[1][942] = 16'h0000;
        rom[1][943] = 16'h0000;
        rom[1][944] = 16'h0000;
        rom[1][945] = 16'h0000;
        rom[1][946] = 16'h0000;
        rom[1][947] = 16'h0000;
        rom[1][948] = 16'h0000;
        rom[1][949] = 16'h0000;
        rom[1][950] = 16'h0000;
        rom[1][951] = 16'h0000;
        rom[1][952] = 16'h0000;
        rom[1][953] = 16'h0000;
        rom[1][954] = 16'h0000;
        rom[1][955] = 16'h0000;
        rom[1][956] = 16'h0000;
        rom[1][957] = 16'h0000;
        rom[1][958] = 16'h0000;
        rom[1][959] = 16'h0000;
        rom[1][960] = 16'h0000;
        rom[1][961] = 16'h0000;
        rom[1][962] = 16'h0000;
        rom[1][963] = 16'h0000;
        rom[1][964] = 16'h0000;
        rom[1][965] = 16'h0000;
        rom[1][966] = 16'h0000;
        rom[1][967] = 16'h0000;
        rom[1][968] = 16'h0000;
        rom[1][969] = 16'h0000;
        rom[1][970] = 16'h0000;
        rom[1][971] = 16'h0000;
        rom[1][972] = 16'h0000;
        rom[1][973] = 16'h0000;
        rom[1][974] = 16'h0000;
        rom[1][975] = 16'h0000;
        rom[1][976] = 16'h0000;
        rom[1][977] = 16'h0000;
        rom[1][978] = 16'h0000;
        rom[1][979] = 16'h0000;
        rom[1][980] = 16'h0104;
        rom[1][981] = 16'h00E7;
        rom[1][982] = 16'h0090;
        rom[1][983] = 16'h00B4;
        rom[1][984] = 16'h00AD;
        rom[1][985] = 16'h00F5;
        rom[1][986] = 16'h00EE;
        rom[1][987] = 16'h00AD;
        rom[1][988] = 16'h0082;
        rom[1][989] = 16'h0048;
        rom[1][990] = 16'h0089;
        rom[1][991] = 16'h00D1;
        rom[1][992] = 16'h00E0;
        rom[1][993] = 16'h0121;
        rom[1][994] = 16'h010B;
        rom[1][995] = 16'h0073;
        rom[1][996] = 16'hFFCD;
        rom[1][997] = 16'h002B;
        rom[1][998] = 16'h00C3;
        rom[1][999] = 16'h00E7;
        rom[1][1000] = 16'h00CA;
        rom[1][1001] = 16'h00C3;
        rom[1][1002] = 16'h00BC;
        rom[1][1003] = 16'h00D9;
        rom[1][1004] = 16'h00FD;
        rom[1][1005] = 16'h0104;
        rom[1][1006] = 16'h007B;
        rom[1][1007] = 16'h0033;
        rom[1][1008] = 16'h003A;
        rom[1][1009] = 16'h0057;
        rom[1][1010] = 16'h00CA;
        rom[1][1011] = 16'h0136;
        rom[1][1012] = 16'h0000;
        rom[1][1013] = 16'h0000;
        rom[1][1014] = 16'h0000;
        rom[1][1015] = 16'h0000;
        rom[1][1016] = 16'h0000;
        rom[1][1017] = 16'h0000;
        rom[1][1018] = 16'h0000;
        rom[1][1019] = 16'h0000;
        rom[1][1020] = 16'h0000;
        rom[1][1021] = 16'h0000;
        rom[1][1022] = 16'h0000;
        rom[1][1023] = 16'h0000;
        rom[1][1024] = 16'h0000;
        rom[1][1025] = 16'h0000;
        rom[1][1026] = 16'h0000;
        rom[1][1027] = 16'h0000;
        rom[1][1028] = 16'h0000;
        rom[1][1029] = 16'h0000;
        rom[1][1030] = 16'h0000;
        rom[1][1031] = 16'h0000;
        rom[1][1032] = 16'h0000;
        rom[1][1033] = 16'h0000;
        rom[1][1034] = 16'h0000;
        rom[1][1035] = 16'h0000;
        rom[1][1036] = 16'h0000;
        rom[1][1037] = 16'h0000;
        rom[1][1038] = 16'h0000;
        rom[1][1039] = 16'h0000;
        rom[1][1040] = 16'h0000;
        rom[1][1041] = 16'h0000;
        rom[1][1042] = 16'h0000;
        rom[1][1043] = 16'h0000;
        rom[1][1044] = 16'h0000;
        rom[1][1045] = 16'h0000;
        rom[1][1046] = 16'h0000;
        rom[1][1047] = 16'h0000;
        rom[1][1048] = 16'h0000;
        rom[1][1049] = 16'h0000;
        rom[1][1050] = 16'h0000;
        rom[1][1051] = 16'h0000;
        rom[1][1052] = 16'h0000;
        rom[1][1053] = 16'h0000;
        rom[1][1054] = 16'h0000;
        rom[1][1055] = 16'h0000;
        rom[1][1056] = 16'h0000;
        rom[1][1057] = 16'h0000;
        rom[1][1058] = 16'h0000;
        rom[1][1059] = 16'h0000;
        rom[1][1060] = 16'h0000;
        rom[1][1061] = 16'h0000;
        rom[1][1062] = 16'h0000;
        rom[1][1063] = 16'h0000;
        rom[1][1064] = 16'h0000;
        rom[1][1065] = 16'h0000;
        rom[1][1066] = 16'h0000;
        rom[1][1067] = 16'h0000;
        rom[1][1068] = 16'h0000;
        rom[1][1069] = 16'h0000;
        rom[1][1070] = 16'h0000;
        rom[1][1071] = 16'h0000;
        rom[1][1072] = 16'h0000;
        rom[1][1073] = 16'h0000;
        rom[1][1074] = 16'h0000;
        rom[1][1075] = 16'h0000;
        rom[1][1076] = 16'h0000;
        rom[1][1077] = 16'h0000;
        rom[1][1078] = 16'h00C3;
        rom[1][1079] = 16'h013E;
        rom[1][1080] = 16'h0169;
        rom[1][1081] = 16'h0136;
        rom[1][1082] = 16'h00F5;
        rom[1][1083] = 16'h00B4;
        rom[1][1084] = 16'hFF27;
        rom[1][1085] = 16'hFE56;
        rom[1][1086] = 16'hFDC6;
        rom[1][1087] = 16'hFDC6;
        rom[1][1088] = 16'hFE0E;
        rom[1][1089] = 16'hFE39;
        rom[1][1090] = 16'hFEFC;
        rom[1][1091] = 16'hFFB8;
        rom[1][1092] = 16'h000E;
        rom[1][1093] = 16'h0000;
        rom[1][1094] = 16'h0024;
        rom[1][1095] = 16'h00EE;
        rom[1][1096] = 16'h018D;
        rom[1][1097] = 16'h0119;
        rom[1][1098] = 16'h00E0;
        rom[1][1099] = 16'h0145;
        rom[1][1100] = 16'h0136;
        rom[1][1101] = 16'h00FD;
        rom[1][1102] = 16'h0119;
        rom[1][1103] = 16'h0119;
        rom[1][1104] = 16'h0104;
        rom[1][1105] = 16'h00EE;
        rom[1][1106] = 16'h00EE;
        rom[1][1107] = 16'h00D9;
        rom[1][1108] = 16'h0112;
        rom[1][1109] = 16'h015A;
        rom[1][1110] = 16'h0000;
        rom[1][1111] = 16'h0000;
        rom[1][1112] = 16'h0000;
        rom[1][1113] = 16'h0000;
        rom[1][1114] = 16'h0000;
        rom[1][1115] = 16'h0000;
        rom[1][1116] = 16'h0000;
        rom[1][1117] = 16'h0000;
        rom[1][1118] = 16'h0000;
        rom[1][1119] = 16'h0000;
        rom[1][1120] = 16'h0000;
        rom[1][1121] = 16'h0000;
        rom[1][1122] = 16'h0000;
        rom[1][1123] = 16'h0000;
        rom[1][1124] = 16'h0000;
        rom[1][1125] = 16'h0000;
        rom[1][1126] = 16'h0000;
        rom[1][1127] = 16'h0000;
        rom[1][1128] = 16'h0000;
        rom[1][1129] = 16'h0000;
        rom[1][1130] = 16'h0000;
        rom[1][1131] = 16'h0000;
        rom[1][1132] = 16'h0000;
        rom[1][1133] = 16'h0000;
        rom[1][1134] = 16'h0000;
        rom[1][1135] = 16'h0000;
        rom[1][1136] = 16'h0000;
        rom[1][1137] = 16'h0000;
        rom[1][1138] = 16'h0000;
        rom[1][1139] = 16'h0000;
        rom[1][1140] = 16'h0000;
        rom[1][1141] = 16'h0000;
        rom[1][1142] = 16'h0000;
        rom[1][1143] = 16'h0000;
        rom[1][1144] = 16'h0000;
        rom[1][1145] = 16'h0000;
        rom[1][1146] = 16'h0000;
        rom[1][1147] = 16'h0000;
        rom[1][1148] = 16'h0000;
        rom[1][1149] = 16'h0000;
        rom[1][1150] = 16'h0000;
        rom[1][1151] = 16'h0000;
        rom[1][1152] = 16'h0000;
        rom[1][1153] = 16'h0000;
        rom[1][1154] = 16'h0000;
        rom[1][1155] = 16'h0000;
        rom[1][1156] = 16'h0000;
        rom[1][1157] = 16'h0000;
        rom[1][1158] = 16'h0000;
        rom[1][1159] = 16'h0000;
        rom[1][1160] = 16'h0000;
        rom[1][1161] = 16'h0000;
        rom[1][1162] = 16'h0000;
        rom[1][1163] = 16'h0000;
        rom[1][1164] = 16'h0000;
        rom[1][1165] = 16'h0000;
        rom[1][1166] = 16'h0000;
        rom[1][1167] = 16'h0000;
        rom[1][1168] = 16'h0000;
        rom[1][1169] = 16'h0000;
        rom[1][1170] = 16'h0000;
        rom[1][1171] = 16'h0000;
        rom[1][1172] = 16'h0000;
        rom[1][1173] = 16'h0000;
        rom[1][1174] = 16'h0000;
        rom[1][1175] = 16'h0000;
        rom[1][1176] = 16'h00B4;
        rom[1][1177] = 16'h00FD;
        rom[1][1178] = 16'h010B;
        rom[1][1179] = 16'h00B4;
        rom[1][1180] = 16'h00AD;
        rom[1][1181] = 16'h0048;
        rom[1][1182] = 16'h0177;
        rom[1][1183] = 16'h0177;
        rom[1][1184] = 16'h0194;
        rom[1][1185] = 16'h013E;
        rom[1][1186] = 16'h00FD;
        rom[1][1187] = 16'h00F5;
        rom[1][1188] = 16'h0128;
        rom[1][1189] = 16'h01CE;
        rom[1][1190] = 16'h01EB;
        rom[1][1191] = 16'h01A3;
        rom[1][1192] = 16'h0112;
        rom[1][1193] = 16'h013E;
        rom[1][1194] = 16'h00FD;
        rom[1][1195] = 16'h0065;
        rom[1][1196] = 16'h007B;
        rom[1][1197] = 16'h0073;
        rom[1][1198] = 16'h00D1;
        rom[1][1199] = 16'h0104;
        rom[1][1200] = 16'h00C3;
        rom[1][1201] = 16'h009F;
        rom[1][1202] = 16'h0082;
        rom[1][1203] = 16'h00EE;
        rom[1][1204] = 16'h0089;
        rom[1][1205] = 16'h0024;
        rom[1][1206] = 16'h004F;
        rom[1][1207] = 16'h006C;
        rom[1][1208] = 16'h0000;
        rom[1][1209] = 16'h0000;
        rom[1][1210] = 16'h0000;
        rom[1][1211] = 16'h0000;
        rom[1][1212] = 16'h0000;
        rom[1][1213] = 16'h0000;
        rom[1][1214] = 16'h0000;
        rom[1][1215] = 16'h0000;
        rom[1][1216] = 16'h0000;
        rom[1][1217] = 16'h0000;
        rom[1][1218] = 16'h0000;
        rom[1][1219] = 16'h0000;
        rom[1][1220] = 16'h0000;
        rom[1][1221] = 16'h0000;
        rom[1][1222] = 16'h0000;
        rom[1][1223] = 16'h0000;
        rom[1][1224] = 16'h0000;
        rom[1][1225] = 16'h0000;
        rom[1][1226] = 16'h0000;
        rom[1][1227] = 16'h0000;
        rom[1][1228] = 16'h0000;
        rom[1][1229] = 16'h0000;
        rom[1][1230] = 16'h0000;
        rom[1][1231] = 16'h0000;
        rom[1][1232] = 16'h0000;
        rom[1][1233] = 16'h0000;
        rom[1][1234] = 16'h0000;
        rom[1][1235] = 16'h0000;
        rom[1][1236] = 16'h0000;
        rom[1][1237] = 16'h0000;
        rom[1][1238] = 16'h0000;
        rom[1][1239] = 16'h0000;
        rom[1][1240] = 16'h0000;
        rom[1][1241] = 16'h0000;
        rom[1][1242] = 16'h0000;
        rom[1][1243] = 16'h0000;
        rom[1][1244] = 16'h0000;
        rom[1][1245] = 16'h0000;
        rom[1][1246] = 16'h0000;
        rom[1][1247] = 16'h0000;
        rom[1][1248] = 16'h0000;
        rom[1][1249] = 16'h0000;
        rom[1][1250] = 16'h0000;
        rom[1][1251] = 16'h0000;
        rom[1][1252] = 16'h0000;
        rom[1][1253] = 16'h0000;
        rom[1][1254] = 16'h0000;
        rom[1][1255] = 16'h0000;
        rom[1][1256] = 16'h0000;
        rom[1][1257] = 16'h0000;
        rom[1][1258] = 16'h0000;
        rom[1][1259] = 16'h0000;
        rom[1][1260] = 16'h0000;
        rom[1][1261] = 16'h0000;
        rom[1][1262] = 16'h0000;
        rom[1][1263] = 16'h0000;
        rom[1][1264] = 16'h0000;
        rom[1][1265] = 16'h0000;
        rom[1][1266] = 16'h0000;
        rom[1][1267] = 16'h0000;
        rom[1][1268] = 16'h0000;
        rom[1][1269] = 16'h0000;
        rom[1][1270] = 16'h0000;
        rom[1][1271] = 16'h0000;
        rom[1][1272] = 16'h0000;
        rom[1][1273] = 16'h0000;
        rom[2][0] = 16'hFFB1;
        rom[2][1] = 16'hFF85;
        rom[2][2] = 16'hFF77;
        rom[2][3] = 16'hFF68;
        rom[2][4] = 16'hFF5A;
        rom[2][5] = 16'hFF44;
        rom[2][6] = 16'hFFA9;
        rom[2][7] = 16'h002B;
        rom[2][8] = 16'h0082;
        rom[2][9] = 16'h00FD;
        rom[2][10] = 16'h0169;
        rom[2][11] = 16'h018D;
        rom[2][12] = 16'h018D;
        rom[2][13] = 16'h0177;
        rom[2][14] = 16'h0121;
        rom[2][15] = 16'h00BC;
        rom[2][16] = 16'h00D9;
        rom[2][17] = 16'h0170;
        rom[2][18] = 16'h017F;
        rom[2][19] = 16'h0136;
        rom[2][20] = 16'h00FD;
        rom[2][21] = 16'h00C3;
        rom[2][22] = 16'h00AD;
        rom[2][23] = 16'h006C;
        rom[2][24] = 16'hFFBF;
        rom[2][25] = 16'hFF36;
        rom[2][26] = 16'hFF7E;
        rom[2][27] = 16'hFFDC;
        rom[2][28] = 16'hFFD5;
        rom[2][29] = 16'hFFB1;
        rom[2][30] = 16'hFFBF;
        rom[2][31] = 16'hFFC6;
        rom[2][32] = 16'h0000;
        rom[2][33] = 16'h0000;
        rom[2][34] = 16'h0000;
        rom[2][35] = 16'h0000;
        rom[2][36] = 16'h0000;
        rom[2][37] = 16'h0000;
        rom[2][38] = 16'h0000;
        rom[2][39] = 16'h0000;
        rom[2][40] = 16'h0000;
        rom[2][41] = 16'h0000;
        rom[2][42] = 16'h0000;
        rom[2][43] = 16'h0000;
        rom[2][44] = 16'h0000;
        rom[2][45] = 16'h0000;
        rom[2][46] = 16'h0000;
        rom[2][47] = 16'h0000;
        rom[2][48] = 16'h0000;
        rom[2][49] = 16'h0000;
        rom[2][50] = 16'h0000;
        rom[2][51] = 16'h0000;
        rom[2][52] = 16'h0000;
        rom[2][53] = 16'h0000;
        rom[2][54] = 16'h0000;
        rom[2][55] = 16'h0000;
        rom[2][56] = 16'h0000;
        rom[2][57] = 16'h0000;
        rom[2][58] = 16'h0000;
        rom[2][59] = 16'h0000;
        rom[2][60] = 16'h0000;
        rom[2][61] = 16'h0000;
        rom[2][62] = 16'h0000;
        rom[2][63] = 16'h0000;
        rom[2][64] = 16'h0000;
        rom[2][65] = 16'h0000;
        rom[2][66] = 16'h0000;
        rom[2][67] = 16'h0000;
        rom[2][68] = 16'h0000;
        rom[2][69] = 16'h0000;
        rom[2][70] = 16'h0000;
        rom[2][71] = 16'h0000;
        rom[2][72] = 16'h0000;
        rom[2][73] = 16'h0000;
        rom[2][74] = 16'h0000;
        rom[2][75] = 16'h0000;
        rom[2][76] = 16'h0000;
        rom[2][77] = 16'h0000;
        rom[2][78] = 16'h0000;
        rom[2][79] = 16'h0000;
        rom[2][80] = 16'h0000;
        rom[2][81] = 16'h0000;
        rom[2][82] = 16'h0000;
        rom[2][83] = 16'h0000;
        rom[2][84] = 16'h0000;
        rom[2][85] = 16'h0000;
        rom[2][86] = 16'h0000;
        rom[2][87] = 16'h0000;
        rom[2][88] = 16'h0000;
        rom[2][89] = 16'h0000;
        rom[2][90] = 16'h0000;
        rom[2][91] = 16'h0000;
        rom[2][92] = 16'h0000;
        rom[2][93] = 16'h0000;
        rom[2][94] = 16'h0000;
        rom[2][95] = 16'h0000;
        rom[2][96] = 16'h0000;
        rom[2][97] = 16'h0000;
        rom[2][98] = 16'hFF0B;
        rom[2][99] = 16'hFF03;
        rom[2][100] = 16'hFF03;
        rom[2][101] = 16'hFF03;
        rom[2][102] = 16'hFF03;
        rom[2][103] = 16'hFEF5;
        rom[2][104] = 16'hFE32;
        rom[2][105] = 16'hFD6F;
        rom[2][106] = 16'hFD6F;
        rom[2][107] = 16'hFECA;
        rom[2][108] = 16'h0041;
        rom[2][109] = 16'h00C3;
        rom[2][110] = 16'h00D1;
        rom[2][111] = 16'h00D9;
        rom[2][112] = 16'h0121;
        rom[2][113] = 16'h0169;
        rom[2][114] = 16'h00E0;
        rom[2][115] = 16'h005E;
        rom[2][116] = 16'h0048;
        rom[2][117] = 16'h0090;
        rom[2][118] = 16'h00CA;
        rom[2][119] = 16'h00D1;
        rom[2][120] = 16'h0145;
        rom[2][121] = 16'h012F;
        rom[2][122] = 16'h0033;
        rom[2][123] = 16'hFF27;
        rom[2][124] = 16'hFF94;
        rom[2][125] = 16'hFFF9;
        rom[2][126] = 16'hFFDC;
        rom[2][127] = 16'hFF44;
        rom[2][128] = 16'hFEEE;
        rom[2][129] = 16'hFEC2;
        rom[2][130] = 16'h0000;
        rom[2][131] = 16'h0000;
        rom[2][132] = 16'h0000;
        rom[2][133] = 16'h0000;
        rom[2][134] = 16'h0000;
        rom[2][135] = 16'h0000;
        rom[2][136] = 16'h0000;
        rom[2][137] = 16'h0000;
        rom[2][138] = 16'h0000;
        rom[2][139] = 16'h0000;
        rom[2][140] = 16'h0000;
        rom[2][141] = 16'h0000;
        rom[2][142] = 16'h0000;
        rom[2][143] = 16'h0000;
        rom[2][144] = 16'h0000;
        rom[2][145] = 16'h0000;
        rom[2][146] = 16'h0000;
        rom[2][147] = 16'h0000;
        rom[2][148] = 16'h0000;
        rom[2][149] = 16'h0000;
        rom[2][150] = 16'h0000;
        rom[2][151] = 16'h0000;
        rom[2][152] = 16'h0000;
        rom[2][153] = 16'h0000;
        rom[2][154] = 16'h0000;
        rom[2][155] = 16'h0000;
        rom[2][156] = 16'h0000;
        rom[2][157] = 16'h0000;
        rom[2][158] = 16'h0000;
        rom[2][159] = 16'h0000;
        rom[2][160] = 16'h0000;
        rom[2][161] = 16'h0000;
        rom[2][162] = 16'h0000;
        rom[2][163] = 16'h0000;
        rom[2][164] = 16'h0000;
        rom[2][165] = 16'h0000;
        rom[2][166] = 16'h0000;
        rom[2][167] = 16'h0000;
        rom[2][168] = 16'h0000;
        rom[2][169] = 16'h0000;
        rom[2][170] = 16'h0000;
        rom[2][171] = 16'h0000;
        rom[2][172] = 16'h0000;
        rom[2][173] = 16'h0000;
        rom[2][174] = 16'h0000;
        rom[2][175] = 16'h0000;
        rom[2][176] = 16'h0000;
        rom[2][177] = 16'h0000;
        rom[2][178] = 16'h0000;
        rom[2][179] = 16'h0000;
        rom[2][180] = 16'h0000;
        rom[2][181] = 16'h0000;
        rom[2][182] = 16'h0000;
        rom[2][183] = 16'h0000;
        rom[2][184] = 16'h0000;
        rom[2][185] = 16'h0000;
        rom[2][186] = 16'h0000;
        rom[2][187] = 16'h0000;
        rom[2][188] = 16'h0000;
        rom[2][189] = 16'h0000;
        rom[2][190] = 16'h0000;
        rom[2][191] = 16'h0000;
        rom[2][192] = 16'h0000;
        rom[2][193] = 16'h0000;
        rom[2][194] = 16'h0000;
        rom[2][195] = 16'h0000;
        rom[2][196] = 16'hFFA2;
        rom[2][197] = 16'hFFB8;
        rom[2][198] = 16'hFFB8;
        rom[2][199] = 16'hFFC6;
        rom[2][200] = 16'hFFCD;
        rom[2][201] = 16'hFFE3;
        rom[2][202] = 16'hFEC2;
        rom[2][203] = 16'hFDD4;
        rom[2][204] = 16'hFD8C;
        rom[2][205] = 16'hFEDF;
        rom[2][206] = 16'hFFEA;
        rom[2][207] = 16'hFFBF;
        rom[2][208] = 16'hFF85;
        rom[2][209] = 16'hFF70;
        rom[2][210] = 16'hFF68;
        rom[2][211] = 16'h0007;
        rom[2][212] = 16'h00BC;
        rom[2][213] = 16'h0073;
        rom[2][214] = 16'h0024;
        rom[2][215] = 16'hFFA9;
        rom[2][216] = 16'hFF36;
        rom[2][217] = 16'hFF2F;
        rom[2][218] = 16'hFEE7;
        rom[2][219] = 16'hFEEE;
        rom[2][220] = 16'hFFBF;
        rom[2][221] = 16'h0041;
        rom[2][222] = 16'h0073;
        rom[2][223] = 16'h003A;
        rom[2][224] = 16'h0065;
        rom[2][225] = 16'h005E;
        rom[2][226] = 16'hFFDC;
        rom[2][227] = 16'hFF8D;
        rom[2][228] = 16'h0000;
        rom[2][229] = 16'h0000;
        rom[2][230] = 16'h0000;
        rom[2][231] = 16'h0000;
        rom[2][232] = 16'h0000;
        rom[2][233] = 16'h0000;
        rom[2][234] = 16'h0000;
        rom[2][235] = 16'h0000;
        rom[2][236] = 16'h0000;
        rom[2][237] = 16'h0000;
        rom[2][238] = 16'h0000;
        rom[2][239] = 16'h0000;
        rom[2][240] = 16'h0000;
        rom[2][241] = 16'h0000;
        rom[2][242] = 16'h0000;
        rom[2][243] = 16'h0000;
        rom[2][244] = 16'h0000;
        rom[2][245] = 16'h0000;
        rom[2][246] = 16'h0000;
        rom[2][247] = 16'h0000;
        rom[2][248] = 16'h0000;
        rom[2][249] = 16'h0000;
        rom[2][250] = 16'h0000;
        rom[2][251] = 16'h0000;
        rom[2][252] = 16'h0000;
        rom[2][253] = 16'h0000;
        rom[2][254] = 16'h0000;
        rom[2][255] = 16'h0000;
        rom[2][256] = 16'h0000;
        rom[2][257] = 16'h0000;
        rom[2][258] = 16'h0000;
        rom[2][259] = 16'h0000;
        rom[2][260] = 16'h0000;
        rom[2][261] = 16'h0000;
        rom[2][262] = 16'h0000;
        rom[2][263] = 16'h0000;
        rom[2][264] = 16'h0000;
        rom[2][265] = 16'h0000;
        rom[2][266] = 16'h0000;
        rom[2][267] = 16'h0000;
        rom[2][268] = 16'h0000;
        rom[2][269] = 16'h0000;
        rom[2][270] = 16'h0000;
        rom[2][271] = 16'h0000;
        rom[2][272] = 16'h0000;
        rom[2][273] = 16'h0000;
        rom[2][274] = 16'h0000;
        rom[2][275] = 16'h0000;
        rom[2][276] = 16'h0000;
        rom[2][277] = 16'h0000;
        rom[2][278] = 16'h0000;
        rom[2][279] = 16'h0000;
        rom[2][280] = 16'h0000;
        rom[2][281] = 16'h0000;
        rom[2][282] = 16'h0000;
        rom[2][283] = 16'h0000;
        rom[2][284] = 16'h0000;
        rom[2][285] = 16'h0000;
        rom[2][286] = 16'h0000;
        rom[2][287] = 16'h0000;
        rom[2][288] = 16'h0000;
        rom[2][289] = 16'h0000;
        rom[2][290] = 16'h0000;
        rom[2][291] = 16'h0000;
        rom[2][292] = 16'h0000;
        rom[2][293] = 16'h0000;
        rom[2][294] = 16'hFF70;
        rom[2][295] = 16'hFF77;
        rom[2][296] = 16'hFF77;
        rom[2][297] = 16'hFF77;
        rom[2][298] = 16'hFF77;
        rom[2][299] = 16'hFF77;
        rom[2][300] = 16'h0089;
        rom[2][301] = 16'h00D9;
        rom[2][302] = 16'h0065;
        rom[2][303] = 16'h0082;
        rom[2][304] = 16'h0007;
        rom[2][305] = 16'hFFF9;
        rom[2][306] = 16'hFFEA;
        rom[2][307] = 16'h0000;
        rom[2][308] = 16'h0007;
        rom[2][309] = 16'hFF9B;
        rom[2][310] = 16'h0057;
        rom[2][311] = 16'h0000;
        rom[2][312] = 16'h0000;
        rom[2][313] = 16'h001D;
        rom[2][314] = 16'hFFDC;
        rom[2][315] = 16'hFFC6;
        rom[2][316] = 16'hFEEE;
        rom[2][317] = 16'hFEDF;
        rom[2][318] = 16'hFF19;
        rom[2][319] = 16'hFFE3;
        rom[2][320] = 16'hFFCD;
        rom[2][321] = 16'hFFCD;
        rom[2][322] = 16'h000E;
        rom[2][323] = 16'h0048;
        rom[2][324] = 16'h0016;
        rom[2][325] = 16'hFFC6;
        rom[2][326] = 16'h0000;
        rom[2][327] = 16'h0000;
        rom[2][328] = 16'h0000;
        rom[2][329] = 16'h0000;
        rom[2][330] = 16'h0000;
        rom[2][331] = 16'h0000;
        rom[2][332] = 16'h0000;
        rom[2][333] = 16'h0000;
        rom[2][334] = 16'h0000;
        rom[2][335] = 16'h0000;
        rom[2][336] = 16'h0000;
        rom[2][337] = 16'h0000;
        rom[2][338] = 16'h0000;
        rom[2][339] = 16'h0000;
        rom[2][340] = 16'h0000;
        rom[2][341] = 16'h0000;
        rom[2][342] = 16'h0000;
        rom[2][343] = 16'h0000;
        rom[2][344] = 16'h0000;
        rom[2][345] = 16'h0000;
        rom[2][346] = 16'h0000;
        rom[2][347] = 16'h0000;
        rom[2][348] = 16'h0000;
        rom[2][349] = 16'h0000;
        rom[2][350] = 16'h0000;
        rom[2][351] = 16'h0000;
        rom[2][352] = 16'h0000;
        rom[2][353] = 16'h0000;
        rom[2][354] = 16'h0000;
        rom[2][355] = 16'h0000;
        rom[2][356] = 16'h0000;
        rom[2][357] = 16'h0000;
        rom[2][358] = 16'h0000;
        rom[2][359] = 16'h0000;
        rom[2][360] = 16'h0000;
        rom[2][361] = 16'h0000;
        rom[2][362] = 16'h0000;
        rom[2][363] = 16'h0000;
        rom[2][364] = 16'h0000;
        rom[2][365] = 16'h0000;
        rom[2][366] = 16'h0000;
        rom[2][367] = 16'h0000;
        rom[2][368] = 16'h0000;
        rom[2][369] = 16'h0000;
        rom[2][370] = 16'h0000;
        rom[2][371] = 16'h0000;
        rom[2][372] = 16'h0000;
        rom[2][373] = 16'h0000;
        rom[2][374] = 16'h0000;
        rom[2][375] = 16'h0000;
        rom[2][376] = 16'h0000;
        rom[2][377] = 16'h0000;
        rom[2][378] = 16'h0000;
        rom[2][379] = 16'h0000;
        rom[2][380] = 16'h0000;
        rom[2][381] = 16'h0000;
        rom[2][382] = 16'h0000;
        rom[2][383] = 16'h0000;
        rom[2][384] = 16'h0000;
        rom[2][385] = 16'h0000;
        rom[2][386] = 16'h0000;
        rom[2][387] = 16'h0000;
        rom[2][388] = 16'h0000;
        rom[2][389] = 16'h0000;
        rom[2][390] = 16'h0000;
        rom[2][391] = 16'h0000;
        rom[2][392] = 16'hFFC6;
        rom[2][393] = 16'hFFE3;
        rom[2][394] = 16'hFFEA;
        rom[2][395] = 16'hFFF9;
        rom[2][396] = 16'h0007;
        rom[2][397] = 16'h0016;
        rom[2][398] = 16'h0098;
        rom[2][399] = 16'h00BC;
        rom[2][400] = 16'hFFB8;
        rom[2][401] = 16'hFF20;
        rom[2][402] = 16'hFE15;
        rom[2][403] = 16'hFDB7;
        rom[2][404] = 16'hFDCD;
        rom[2][405] = 16'hFE6C;
        rom[2][406] = 16'hFF68;
        rom[2][407] = 16'hFFBF;
        rom[2][408] = 16'hFEAD;
        rom[2][409] = 16'hFEEE;
        rom[2][410] = 16'hFEC2;
        rom[2][411] = 16'hFDF1;
        rom[2][412] = 16'hFE41;
        rom[2][413] = 16'hFF5A;
        rom[2][414] = 16'h0065;
        rom[2][415] = 16'h0082;
        rom[2][416] = 16'h0082;
        rom[2][417] = 16'h0073;
        rom[2][418] = 16'hFFEA;
        rom[2][419] = 16'hFF53;
        rom[2][420] = 16'hFF53;
        rom[2][421] = 16'hFFA2;
        rom[2][422] = 16'hFF5A;
        rom[2][423] = 16'hFF53;
        rom[2][424] = 16'h0000;
        rom[2][425] = 16'h0000;
        rom[2][426] = 16'h0000;
        rom[2][427] = 16'h0000;
        rom[2][428] = 16'h0000;
        rom[2][429] = 16'h0000;
        rom[2][430] = 16'h0000;
        rom[2][431] = 16'h0000;
        rom[2][432] = 16'h0000;
        rom[2][433] = 16'h0000;
        rom[2][434] = 16'h0000;
        rom[2][435] = 16'h0000;
        rom[2][436] = 16'h0000;
        rom[2][437] = 16'h0000;
        rom[2][438] = 16'h0000;
        rom[2][439] = 16'h0000;
        rom[2][440] = 16'h0000;
        rom[2][441] = 16'h0000;
        rom[2][442] = 16'h0000;
        rom[2][443] = 16'h0000;
        rom[2][444] = 16'h0000;
        rom[2][445] = 16'h0000;
        rom[2][446] = 16'h0000;
        rom[2][447] = 16'h0000;
        rom[2][448] = 16'h0000;
        rom[2][449] = 16'h0000;
        rom[2][450] = 16'h0000;
        rom[2][451] = 16'h0000;
        rom[2][452] = 16'h0000;
        rom[2][453] = 16'h0000;
        rom[2][454] = 16'h0000;
        rom[2][455] = 16'h0000;
        rom[2][456] = 16'h0000;
        rom[2][457] = 16'h0000;
        rom[2][458] = 16'h0000;
        rom[2][459] = 16'h0000;
        rom[2][460] = 16'h0000;
        rom[2][461] = 16'h0000;
        rom[2][462] = 16'h0000;
        rom[2][463] = 16'h0000;
        rom[2][464] = 16'h0000;
        rom[2][465] = 16'h0000;
        rom[2][466] = 16'h0000;
        rom[2][467] = 16'h0000;
        rom[2][468] = 16'h0000;
        rom[2][469] = 16'h0000;
        rom[2][470] = 16'h0000;
        rom[2][471] = 16'h0000;
        rom[2][472] = 16'h0000;
        rom[2][473] = 16'h0000;
        rom[2][474] = 16'h0000;
        rom[2][475] = 16'h0000;
        rom[2][476] = 16'h0000;
        rom[2][477] = 16'h0000;
        rom[2][478] = 16'h0000;
        rom[2][479] = 16'h0000;
        rom[2][480] = 16'h0000;
        rom[2][481] = 16'h0000;
        rom[2][482] = 16'h0000;
        rom[2][483] = 16'h0000;
        rom[2][484] = 16'h0000;
        rom[2][485] = 16'h0000;
        rom[2][486] = 16'h0000;
        rom[2][487] = 16'h0000;
        rom[2][488] = 16'h0000;
        rom[2][489] = 16'h0000;
        rom[2][490] = 16'hFF8D;
        rom[2][491] = 16'hFF94;
        rom[2][492] = 16'hFFA2;
        rom[2][493] = 16'hFFB1;
        rom[2][494] = 16'hFFBF;
        rom[2][495] = 16'hFFCD;
        rom[2][496] = 16'h0082;
        rom[2][497] = 16'h00D9;
        rom[2][498] = 16'hFFCD;
        rom[2][499] = 16'hFF53;
        rom[2][500] = 16'hFF20;
        rom[2][501] = 16'hFEFC;
        rom[2][502] = 16'hFECA;
        rom[2][503] = 16'hFE81;
        rom[2][504] = 16'hFE56;
        rom[2][505] = 16'hFE9E;
        rom[2][506] = 16'hFECA;
        rom[2][507] = 16'hFF70;
        rom[2][508] = 16'hFF70;
        rom[2][509] = 16'hFE9E;
        rom[2][510] = 16'hFDEA;
        rom[2][511] = 16'hFE15;
        rom[2][512] = 16'hFDC6;
        rom[2][513] = 16'hFE32;
        rom[2][514] = 16'hFF20;
        rom[2][515] = 16'hFFEA;
        rom[2][516] = 16'hFEE7;
        rom[2][517] = 16'hFE81;
        rom[2][518] = 16'hFE89;
        rom[2][519] = 16'hFF94;
        rom[2][520] = 16'h0057;
        rom[2][521] = 16'h0082;
        rom[2][522] = 16'h0000;
        rom[2][523] = 16'h0000;
        rom[2][524] = 16'h0000;
        rom[2][525] = 16'h0000;
        rom[2][526] = 16'h0000;
        rom[2][527] = 16'h0000;
        rom[2][528] = 16'h0000;
        rom[2][529] = 16'h0000;
        rom[2][530] = 16'h0000;
        rom[2][531] = 16'h0000;
        rom[2][532] = 16'h0000;
        rom[2][533] = 16'h0000;
        rom[2][534] = 16'h0000;
        rom[2][535] = 16'h0000;
        rom[2][536] = 16'h0000;
        rom[2][537] = 16'h0000;
        rom[2][538] = 16'h0000;
        rom[2][539] = 16'h0000;
        rom[2][540] = 16'h0000;
        rom[2][541] = 16'h0000;
        rom[2][542] = 16'h0000;
        rom[2][543] = 16'h0000;
        rom[2][544] = 16'h0000;
        rom[2][545] = 16'h0000;
        rom[2][546] = 16'h0000;
        rom[2][547] = 16'h0000;
        rom[2][548] = 16'h0000;
        rom[2][549] = 16'h0000;
        rom[2][550] = 16'h0000;
        rom[2][551] = 16'h0000;
        rom[2][552] = 16'h0000;
        rom[2][553] = 16'h0000;
        rom[2][554] = 16'h0000;
        rom[2][555] = 16'h0000;
        rom[2][556] = 16'h0000;
        rom[2][557] = 16'h0000;
        rom[2][558] = 16'h0000;
        rom[2][559] = 16'h0000;
        rom[2][560] = 16'h0000;
        rom[2][561] = 16'h0000;
        rom[2][562] = 16'h0000;
        rom[2][563] = 16'h0000;
        rom[2][564] = 16'h0000;
        rom[2][565] = 16'h0000;
        rom[2][566] = 16'h0000;
        rom[2][567] = 16'h0000;
        rom[2][568] = 16'h0000;
        rom[2][569] = 16'h0000;
        rom[2][570] = 16'h0000;
        rom[2][571] = 16'h0000;
        rom[2][572] = 16'h0000;
        rom[2][573] = 16'h0000;
        rom[2][574] = 16'h0000;
        rom[2][575] = 16'h0000;
        rom[2][576] = 16'h0000;
        rom[2][577] = 16'h0000;
        rom[2][578] = 16'h0000;
        rom[2][579] = 16'h0000;
        rom[2][580] = 16'h0000;
        rom[2][581] = 16'h0000;
        rom[2][582] = 16'h0000;
        rom[2][583] = 16'h0000;
        rom[2][584] = 16'h0000;
        rom[2][585] = 16'h0000;
        rom[2][586] = 16'h0000;
        rom[2][587] = 16'h0000;
        rom[2][588] = 16'h0007;
        rom[2][589] = 16'h001D;
        rom[2][590] = 16'h002B;
        rom[2][591] = 16'h003A;
        rom[2][592] = 16'h0041;
        rom[2][593] = 16'h004F;
        rom[2][594] = 16'hFECA;
        rom[2][595] = 16'hFEFC;
        rom[2][596] = 16'hFF7E;
        rom[2][597] = 16'hFF36;
        rom[2][598] = 16'hFF8D;
        rom[2][599] = 16'h00A6;
        rom[2][600] = 16'h0128;
        rom[2][601] = 16'h00E0;
        rom[2][602] = 16'h00A6;
        rom[2][603] = 16'h009F;
        rom[2][604] = 16'h0048;
        rom[2][605] = 16'hFFCD;
        rom[2][606] = 16'h004F;
        rom[2][607] = 16'h01EB;
        rom[2][608] = 16'h0291;
        rom[2][609] = 16'h0153;
        rom[2][610] = 16'hFF85;
        rom[2][611] = 16'hFED1;
        rom[2][612] = 16'hFE90;
        rom[2][613] = 16'hFFF9;
        rom[2][614] = 16'hFE9E;
        rom[2][615] = 16'hFDB7;
        rom[2][616] = 16'hFDEA;
        rom[2][617] = 16'hFEF5;
        rom[2][618] = 16'hFF68;
        rom[2][619] = 16'hFFB8;
        rom[2][620] = 16'h0000;
        rom[2][621] = 16'h0000;
        rom[2][622] = 16'h0000;
        rom[2][623] = 16'h0000;
        rom[2][624] = 16'h0000;
        rom[2][625] = 16'h0000;
        rom[2][626] = 16'h0000;
        rom[2][627] = 16'h0000;
        rom[2][628] = 16'h0000;
        rom[2][629] = 16'h0000;
        rom[2][630] = 16'h0000;
        rom[2][631] = 16'h0000;
        rom[2][632] = 16'h0000;
        rom[2][633] = 16'h0000;
        rom[2][634] = 16'h0000;
        rom[2][635] = 16'h0000;
        rom[2][636] = 16'h0000;
        rom[2][637] = 16'h0000;
        rom[2][638] = 16'h0000;
        rom[2][639] = 16'h0000;
        rom[2][640] = 16'h0000;
        rom[2][641] = 16'h0000;
        rom[2][642] = 16'h0000;
        rom[2][643] = 16'h0000;
        rom[2][644] = 16'h0000;
        rom[2][645] = 16'h0000;
        rom[2][646] = 16'h0000;
        rom[2][647] = 16'h0000;
        rom[2][648] = 16'h0000;
        rom[2][649] = 16'h0000;
        rom[2][650] = 16'h0000;
        rom[2][651] = 16'h0000;
        rom[2][652] = 16'h0000;
        rom[2][653] = 16'h0000;
        rom[2][654] = 16'h0000;
        rom[2][655] = 16'h0000;
        rom[2][656] = 16'h0000;
        rom[2][657] = 16'h0000;
        rom[2][658] = 16'h0000;
        rom[2][659] = 16'h0000;
        rom[2][660] = 16'h0000;
        rom[2][661] = 16'h0000;
        rom[2][662] = 16'h0000;
        rom[2][663] = 16'h0000;
        rom[2][664] = 16'h0000;
        rom[2][665] = 16'h0000;
        rom[2][666] = 16'h0000;
        rom[2][667] = 16'h0000;
        rom[2][668] = 16'h0000;
        rom[2][669] = 16'h0000;
        rom[2][670] = 16'h0000;
        rom[2][671] = 16'h0000;
        rom[2][672] = 16'h0000;
        rom[2][673] = 16'h0000;
        rom[2][674] = 16'h0000;
        rom[2][675] = 16'h0000;
        rom[2][676] = 16'h0000;
        rom[2][677] = 16'h0000;
        rom[2][678] = 16'h0000;
        rom[2][679] = 16'h0000;
        rom[2][680] = 16'h0000;
        rom[2][681] = 16'h0000;
        rom[2][682] = 16'h0000;
        rom[2][683] = 16'h0000;
        rom[2][684] = 16'h0000;
        rom[2][685] = 16'h0000;
        rom[2][686] = 16'hFFCD;
        rom[2][687] = 16'hFFDC;
        rom[2][688] = 16'hFFEA;
        rom[2][689] = 16'hFFF9;
        rom[2][690] = 16'h0007;
        rom[2][691] = 16'h0016;
        rom[2][692] = 16'hFFB1;
        rom[2][693] = 16'hFFF9;
        rom[2][694] = 16'h0073;
        rom[2][695] = 16'hFFF2;
        rom[2][696] = 16'hFFE3;
        rom[2][697] = 16'hFF85;
        rom[2][698] = 16'hFF20;
        rom[2][699] = 16'hFED1;
        rom[2][700] = 16'hFE24;
        rom[2][701] = 16'hFDDB;
        rom[2][702] = 16'hFEBB;
        rom[2][703] = 16'hFF70;
        rom[2][704] = 16'hFF4C;
        rom[2][705] = 16'hFE97;
        rom[2][706] = 16'hFDF1;
        rom[2][707] = 16'hFD6F;
        rom[2][708] = 16'hFE07;
        rom[2][709] = 16'hFE39;
        rom[2][710] = 16'hFE41;
        rom[2][711] = 16'hFF4C;
        rom[2][712] = 16'hFDE3;
        rom[2][713] = 16'h0362;
        rom[2][714] = 16'h0371;
        rom[2][715] = 16'hFDB7;
        rom[2][716] = 16'hFE89;
        rom[2][717] = 16'hFF53;
        rom[2][718] = 16'h0000;
        rom[2][719] = 16'h0000;
        rom[2][720] = 16'h0000;
        rom[2][721] = 16'h0000;
        rom[2][722] = 16'h0000;
        rom[2][723] = 16'h0000;
        rom[2][724] = 16'h0000;
        rom[2][725] = 16'h0000;
        rom[2][726] = 16'h0000;
        rom[2][727] = 16'h0000;
        rom[2][728] = 16'h0000;
        rom[2][729] = 16'h0000;
        rom[2][730] = 16'h0000;
        rom[2][731] = 16'h0000;
        rom[2][732] = 16'h0000;
        rom[2][733] = 16'h0000;
        rom[2][734] = 16'h0000;
        rom[2][735] = 16'h0000;
        rom[2][736] = 16'h0000;
        rom[2][737] = 16'h0000;
        rom[2][738] = 16'h0000;
        rom[2][739] = 16'h0000;
        rom[2][740] = 16'h0000;
        rom[2][741] = 16'h0000;
        rom[2][742] = 16'h0000;
        rom[2][743] = 16'h0000;
        rom[2][744] = 16'h0000;
        rom[2][745] = 16'h0000;
        rom[2][746] = 16'h0000;
        rom[2][747] = 16'h0000;
        rom[2][748] = 16'h0000;
        rom[2][749] = 16'h0000;
        rom[2][750] = 16'h0000;
        rom[2][751] = 16'h0000;
        rom[2][752] = 16'h0000;
        rom[2][753] = 16'h0000;
        rom[2][754] = 16'h0000;
        rom[2][755] = 16'h0000;
        rom[2][756] = 16'h0000;
        rom[2][757] = 16'h0000;
        rom[2][758] = 16'h0000;
        rom[2][759] = 16'h0000;
        rom[2][760] = 16'h0000;
        rom[2][761] = 16'h0000;
        rom[2][762] = 16'h0000;
        rom[2][763] = 16'h0000;
        rom[2][764] = 16'h0000;
        rom[2][765] = 16'h0000;
        rom[2][766] = 16'h0000;
        rom[2][767] = 16'h0000;
        rom[2][768] = 16'h0000;
        rom[2][769] = 16'h0000;
        rom[2][770] = 16'h0000;
        rom[2][771] = 16'h0000;
        rom[2][772] = 16'h0000;
        rom[2][773] = 16'h0000;
        rom[2][774] = 16'h0000;
        rom[2][775] = 16'h0000;
        rom[2][776] = 16'h0000;
        rom[2][777] = 16'h0000;
        rom[2][778] = 16'h0000;
        rom[2][779] = 16'h0000;
        rom[2][780] = 16'h0000;
        rom[2][781] = 16'h0000;
        rom[2][782] = 16'h0000;
        rom[2][783] = 16'h0000;
        rom[2][784] = 16'h001D;
        rom[2][785] = 16'h0033;
        rom[2][786] = 16'h003A;
        rom[2][787] = 16'h0041;
        rom[2][788] = 16'h0048;
        rom[2][789] = 16'h004F;
        rom[2][790] = 16'h0216;
        rom[2][791] = 16'h00D9;
        rom[2][792] = 16'hFFD5;
        rom[2][793] = 16'hFEBB;
        rom[2][794] = 16'hFE97;
        rom[2][795] = 16'hFE5D;
        rom[2][796] = 16'hFE7A;
        rom[2][797] = 16'hFE5D;
        rom[2][798] = 16'hFE90;
        rom[2][799] = 16'hFF12;
        rom[2][800] = 16'hFF44;
        rom[2][801] = 16'hFF7E;
        rom[2][802] = 16'hFF0B;
        rom[2][803] = 16'hFE24;
        rom[2][804] = 16'hFE24;
        rom[2][805] = 16'hFE0E;
        rom[2][806] = 16'hFDC6;
        rom[2][807] = 16'hFE5D;
        rom[2][808] = 16'hFF36;
        rom[2][809] = 16'hFFB8;
        rom[2][810] = 16'hFF7E;
        rom[2][811] = 16'h003A;
        rom[2][812] = 16'hFFBF;
        rom[2][813] = 16'hFF0B;
        rom[2][814] = 16'hFFBF;
        rom[2][815] = 16'hFFB8;
        rom[2][816] = 16'h0000;
        rom[2][817] = 16'h0000;
        rom[2][818] = 16'h0000;
        rom[2][819] = 16'h0000;
        rom[2][820] = 16'h0000;
        rom[2][821] = 16'h0000;
        rom[2][822] = 16'h0000;
        rom[2][823] = 16'h0000;
        rom[2][824] = 16'h0000;
        rom[2][825] = 16'h0000;
        rom[2][826] = 16'h0000;
        rom[2][827] = 16'h0000;
        rom[2][828] = 16'h0000;
        rom[2][829] = 16'h0000;
        rom[2][830] = 16'h0000;
        rom[2][831] = 16'h0000;
        rom[2][832] = 16'h0000;
        rom[2][833] = 16'h0000;
        rom[2][834] = 16'h0000;
        rom[2][835] = 16'h0000;
        rom[2][836] = 16'h0000;
        rom[2][837] = 16'h0000;
        rom[2][838] = 16'h0000;
        rom[2][839] = 16'h0000;
        rom[2][840] = 16'h0000;
        rom[2][841] = 16'h0000;
        rom[2][842] = 16'h0000;
        rom[2][843] = 16'h0000;
        rom[2][844] = 16'h0000;
        rom[2][845] = 16'h0000;
        rom[2][846] = 16'h0000;
        rom[2][847] = 16'h0000;
        rom[2][848] = 16'h0000;
        rom[2][849] = 16'h0000;
        rom[2][850] = 16'h0000;
        rom[2][851] = 16'h0000;
        rom[2][852] = 16'h0000;
        rom[2][853] = 16'h0000;
        rom[2][854] = 16'h0000;
        rom[2][855] = 16'h0000;
        rom[2][856] = 16'h0000;
        rom[2][857] = 16'h0000;
        rom[2][858] = 16'h0000;
        rom[2][859] = 16'h0000;
        rom[2][860] = 16'h0000;
        rom[2][861] = 16'h0000;
        rom[2][862] = 16'h0000;
        rom[2][863] = 16'h0000;
        rom[2][864] = 16'h0000;
        rom[2][865] = 16'h0000;
        rom[2][866] = 16'h0000;
        rom[2][867] = 16'h0000;
        rom[2][868] = 16'h0000;
        rom[2][869] = 16'h0000;
        rom[2][870] = 16'h0000;
        rom[2][871] = 16'h0000;
        rom[2][872] = 16'h0000;
        rom[2][873] = 16'h0000;
        rom[2][874] = 16'h0000;
        rom[2][875] = 16'h0000;
        rom[2][876] = 16'h0000;
        rom[2][877] = 16'h0000;
        rom[2][878] = 16'h0000;
        rom[2][879] = 16'h0000;
        rom[2][880] = 16'h0000;
        rom[2][881] = 16'h0000;
        rom[2][882] = 16'hFFEA;
        rom[2][883] = 16'hFFF2;
        rom[2][884] = 16'hFFF9;
        rom[2][885] = 16'h0000;
        rom[2][886] = 16'h0007;
        rom[2][887] = 16'h0007;
        rom[2][888] = 16'h0024;
        rom[2][889] = 16'h00C3;
        rom[2][890] = 16'h0119;
        rom[2][891] = 16'h005E;
        rom[2][892] = 16'hFFF2;
        rom[2][893] = 16'hFFF9;
        rom[2][894] = 16'h0090;
        rom[2][895] = 16'hFFE3;
        rom[2][896] = 16'hFF20;
        rom[2][897] = 16'hFE97;
        rom[2][898] = 16'hFF4C;
        rom[2][899] = 16'hFFB1;
        rom[2][900] = 16'h000E;
        rom[2][901] = 16'h00C3;
        rom[2][902] = 16'h0112;
        rom[2][903] = 16'h017F;
        rom[2][904] = 16'h015A;
        rom[2][905] = 16'h00CA;
        rom[2][906] = 16'hFFEA;
        rom[2][907] = 16'hFFDC;
        rom[2][908] = 16'hFFF9;
        rom[2][909] = 16'h004F;
        rom[2][910] = 16'h000E;
        rom[2][911] = 16'hFF0B;
        rom[2][912] = 16'hFFB8;
        rom[2][913] = 16'hFF94;
        rom[2][914] = 16'h0000;
        rom[2][915] = 16'h0000;
        rom[2][916] = 16'h0000;
        rom[2][917] = 16'h0000;
        rom[2][918] = 16'h0000;
        rom[2][919] = 16'h0000;
        rom[2][920] = 16'h0000;
        rom[2][921] = 16'h0000;
        rom[2][922] = 16'h0000;
        rom[2][923] = 16'h0000;
        rom[2][924] = 16'h0000;
        rom[2][925] = 16'h0000;
        rom[2][926] = 16'h0000;
        rom[2][927] = 16'h0000;
        rom[2][928] = 16'h0000;
        rom[2][929] = 16'h0000;
        rom[2][930] = 16'h0000;
        rom[2][931] = 16'h0000;
        rom[2][932] = 16'h0000;
        rom[2][933] = 16'h0000;
        rom[2][934] = 16'h0000;
        rom[2][935] = 16'h0000;
        rom[2][936] = 16'h0000;
        rom[2][937] = 16'h0000;
        rom[2][938] = 16'h0000;
        rom[2][939] = 16'h0000;
        rom[2][940] = 16'h0000;
        rom[2][941] = 16'h0000;
        rom[2][942] = 16'h0000;
        rom[2][943] = 16'h0000;
        rom[2][944] = 16'h0000;
        rom[2][945] = 16'h0000;
        rom[2][946] = 16'h0000;
        rom[2][947] = 16'h0000;
        rom[2][948] = 16'h0000;
        rom[2][949] = 16'h0000;
        rom[2][950] = 16'h0000;
        rom[2][951] = 16'h0000;
        rom[2][952] = 16'h0000;
        rom[2][953] = 16'h0000;
        rom[2][954] = 16'h0000;
        rom[2][955] = 16'h0000;
        rom[2][956] = 16'h0000;
        rom[2][957] = 16'h0000;
        rom[2][958] = 16'h0000;
        rom[2][959] = 16'h0000;
        rom[2][960] = 16'h0000;
        rom[2][961] = 16'h0000;
        rom[2][962] = 16'h0000;
        rom[2][963] = 16'h0000;
        rom[2][964] = 16'h0000;
        rom[2][965] = 16'h0000;
        rom[2][966] = 16'h0000;
        rom[2][967] = 16'h0000;
        rom[2][968] = 16'h0000;
        rom[2][969] = 16'h0000;
        rom[2][970] = 16'h0000;
        rom[2][971] = 16'h0000;
        rom[2][972] = 16'h0000;
        rom[2][973] = 16'h0000;
        rom[2][974] = 16'h0000;
        rom[2][975] = 16'h0000;
        rom[2][976] = 16'h0000;
        rom[2][977] = 16'h0000;
        rom[2][978] = 16'h0000;
        rom[2][979] = 16'h0000;
        rom[2][980] = 16'h0048;
        rom[2][981] = 16'h005E;
        rom[2][982] = 16'h006C;
        rom[2][983] = 16'h006C;
        rom[2][984] = 16'h006C;
        rom[2][985] = 16'h0073;
        rom[2][986] = 16'hFF27;
        rom[2][987] = 16'hFF2F;
        rom[2][988] = 16'hFFE3;
        rom[2][989] = 16'hFF03;
        rom[2][990] = 16'hFEC2;
        rom[2][991] = 16'hFEF5;
        rom[2][992] = 16'hFF20;
        rom[2][993] = 16'hFEDF;
        rom[2][994] = 16'hFE56;
        rom[2][995] = 16'hFD9B;
        rom[2][996] = 16'hFDC6;
        rom[2][997] = 16'hFE65;
        rom[2][998] = 16'hFF27;
        rom[2][999] = 16'hFF94;
        rom[2][1000] = 16'hFF4C;
        rom[2][1001] = 16'hFFF9;
        rom[2][1002] = 16'h015A;
        rom[2][1003] = 16'h0249;
        rom[2][1004] = 16'h00EE;
        rom[2][1005] = 16'h0098;
        rom[2][1006] = 16'hFFC6;
        rom[2][1007] = 16'hFE32;
        rom[2][1008] = 16'hFE73;
        rom[2][1009] = 16'hFFC6;
        rom[2][1010] = 16'h0112;
        rom[2][1011] = 16'h0186;
        rom[2][1012] = 16'h0000;
        rom[2][1013] = 16'h0000;
        rom[2][1014] = 16'h0000;
        rom[2][1015] = 16'h0000;
        rom[2][1016] = 16'h0000;
        rom[2][1017] = 16'h0000;
        rom[2][1018] = 16'h0000;
        rom[2][1019] = 16'h0000;
        rom[2][1020] = 16'h0000;
        rom[2][1021] = 16'h0000;
        rom[2][1022] = 16'h0000;
        rom[2][1023] = 16'h0000;
        rom[2][1024] = 16'h0000;
        rom[2][1025] = 16'h0000;
        rom[2][1026] = 16'h0000;
        rom[2][1027] = 16'h0000;
        rom[2][1028] = 16'h0000;
        rom[2][1029] = 16'h0000;
        rom[2][1030] = 16'h0000;
        rom[2][1031] = 16'h0000;
        rom[2][1032] = 16'h0000;
        rom[2][1033] = 16'h0000;
        rom[2][1034] = 16'h0000;
        rom[2][1035] = 16'h0000;
        rom[2][1036] = 16'h0000;
        rom[2][1037] = 16'h0000;
        rom[2][1038] = 16'h0000;
        rom[2][1039] = 16'h0000;
        rom[2][1040] = 16'h0000;
        rom[2][1041] = 16'h0000;
        rom[2][1042] = 16'h0000;
        rom[2][1043] = 16'h0000;
        rom[2][1044] = 16'h0000;
        rom[2][1045] = 16'h0000;
        rom[2][1046] = 16'h0000;
        rom[2][1047] = 16'h0000;
        rom[2][1048] = 16'h0000;
        rom[2][1049] = 16'h0000;
        rom[2][1050] = 16'h0000;
        rom[2][1051] = 16'h0000;
        rom[2][1052] = 16'h0000;
        rom[2][1053] = 16'h0000;
        rom[2][1054] = 16'h0000;
        rom[2][1055] = 16'h0000;
        rom[2][1056] = 16'h0000;
        rom[2][1057] = 16'h0000;
        rom[2][1058] = 16'h0000;
        rom[2][1059] = 16'h0000;
        rom[2][1060] = 16'h0000;
        rom[2][1061] = 16'h0000;
        rom[2][1062] = 16'h0000;
        rom[2][1063] = 16'h0000;
        rom[2][1064] = 16'h0000;
        rom[2][1065] = 16'h0000;
        rom[2][1066] = 16'h0000;
        rom[2][1067] = 16'h0000;
        rom[2][1068] = 16'h0000;
        rom[2][1069] = 16'h0000;
        rom[2][1070] = 16'h0000;
        rom[2][1071] = 16'h0000;
        rom[2][1072] = 16'h0000;
        rom[2][1073] = 16'h0000;
        rom[2][1074] = 16'h0000;
        rom[2][1075] = 16'h0000;
        rom[2][1076] = 16'h0000;
        rom[2][1077] = 16'h0000;
        rom[2][1078] = 16'hFFF9;
        rom[2][1079] = 16'hFFF9;
        rom[2][1080] = 16'h0000;
        rom[2][1081] = 16'h0007;
        rom[2][1082] = 16'h000E;
        rom[2][1083] = 16'h000E;
        rom[2][1084] = 16'h00E7;
        rom[2][1085] = 16'h0098;
        rom[2][1086] = 16'h009F;
        rom[2][1087] = 16'h0048;
        rom[2][1088] = 16'h00E7;
        rom[2][1089] = 16'h014C;
        rom[2][1090] = 16'h021D;
        rom[2][1091] = 16'h025E;
        rom[2][1092] = 16'h01F9;
        rom[2][1093] = 16'h0104;
        rom[2][1094] = 16'hFFE3;
        rom[2][1095] = 16'h003A;
        rom[2][1096] = 16'h0169;
        rom[2][1097] = 16'h02C3;
        rom[2][1098] = 16'h02E7;
        rom[2][1099] = 16'h0274;
        rom[2][1100] = 16'h0121;
        rom[2][1101] = 16'h0073;
        rom[2][1102] = 16'h0057;
        rom[2][1103] = 16'hFFEA;
        rom[2][1104] = 16'hFF12;
        rom[2][1105] = 16'hFECA;
        rom[2][1106] = 16'hFED1;
        rom[2][1107] = 16'hFF44;
        rom[2][1108] = 16'hFE6C;
        rom[2][1109] = 16'hFE9E;
        rom[2][1110] = 16'h0000;
        rom[2][1111] = 16'h0000;
        rom[2][1112] = 16'h0000;
        rom[2][1113] = 16'h0000;
        rom[2][1114] = 16'h0000;
        rom[2][1115] = 16'h0000;
        rom[2][1116] = 16'h0000;
        rom[2][1117] = 16'h0000;
        rom[2][1118] = 16'h0000;
        rom[2][1119] = 16'h0000;
        rom[2][1120] = 16'h0000;
        rom[2][1121] = 16'h0000;
        rom[2][1122] = 16'h0000;
        rom[2][1123] = 16'h0000;
        rom[2][1124] = 16'h0000;
        rom[2][1125] = 16'h0000;
        rom[2][1126] = 16'h0000;
        rom[2][1127] = 16'h0000;
        rom[2][1128] = 16'h0000;
        rom[2][1129] = 16'h0000;
        rom[2][1130] = 16'h0000;
        rom[2][1131] = 16'h0000;
        rom[2][1132] = 16'h0000;
        rom[2][1133] = 16'h0000;
        rom[2][1134] = 16'h0000;
        rom[2][1135] = 16'h0000;
        rom[2][1136] = 16'h0000;
        rom[2][1137] = 16'h0000;
        rom[2][1138] = 16'h0000;
        rom[2][1139] = 16'h0000;
        rom[2][1140] = 16'h0000;
        rom[2][1141] = 16'h0000;
        rom[2][1142] = 16'h0000;
        rom[2][1143] = 16'h0000;
        rom[2][1144] = 16'h0000;
        rom[2][1145] = 16'h0000;
        rom[2][1146] = 16'h0000;
        rom[2][1147] = 16'h0000;
        rom[2][1148] = 16'h0000;
        rom[2][1149] = 16'h0000;
        rom[2][1150] = 16'h0000;
        rom[2][1151] = 16'h0000;
        rom[2][1152] = 16'h0000;
        rom[2][1153] = 16'h0000;
        rom[2][1154] = 16'h0000;
        rom[2][1155] = 16'h0000;
        rom[2][1156] = 16'h0000;
        rom[2][1157] = 16'h0000;
        rom[2][1158] = 16'h0000;
        rom[2][1159] = 16'h0000;
        rom[2][1160] = 16'h0000;
        rom[2][1161] = 16'h0000;
        rom[2][1162] = 16'h0000;
        rom[2][1163] = 16'h0000;
        rom[2][1164] = 16'h0000;
        rom[2][1165] = 16'h0000;
        rom[2][1166] = 16'h0000;
        rom[2][1167] = 16'h0000;
        rom[2][1168] = 16'h0000;
        rom[2][1169] = 16'h0000;
        rom[2][1170] = 16'h0000;
        rom[2][1171] = 16'h0000;
        rom[2][1172] = 16'h0000;
        rom[2][1173] = 16'h0000;
        rom[2][1174] = 16'h0000;
        rom[2][1175] = 16'h0000;
        rom[2][1176] = 16'h0048;
        rom[2][1177] = 16'h0057;
        rom[2][1178] = 16'h0065;
        rom[2][1179] = 16'h0065;
        rom[2][1180] = 16'h006C;
        rom[2][1181] = 16'h0073;
        rom[2][1182] = 16'hFF9B;
        rom[2][1183] = 16'hFF61;
        rom[2][1184] = 16'hFF68;
        rom[2][1185] = 16'hFEBB;
        rom[2][1186] = 16'h0007;
        rom[2][1187] = 16'h0065;
        rom[2][1188] = 16'h002B;
        rom[2][1189] = 16'hFFF2;
        rom[2][1190] = 16'hFFEA;
        rom[2][1191] = 16'hFFF9;
        rom[2][1192] = 16'hFECA;
        rom[2][1193] = 16'hFF85;
        rom[2][1194] = 16'h0007;
        rom[2][1195] = 16'hFE7A;
        rom[2][1196] = 16'hFD35;
        rom[2][1197] = 16'hFD44;
        rom[2][1198] = 16'hFE7A;
        rom[2][1199] = 16'hFF85;
        rom[2][1200] = 16'h00AD;
        rom[2][1201] = 16'hFFE3;
        rom[2][1202] = 16'hFFD5;
        rom[2][1203] = 16'hFF53;
        rom[2][1204] = 16'hFF3D;
        rom[2][1205] = 16'h0033;
        rom[2][1206] = 16'hFFEA;
        rom[2][1207] = 16'h0016;
        rom[2][1208] = 16'h0000;
        rom[2][1209] = 16'h0000;
        rom[2][1210] = 16'h0000;
        rom[2][1211] = 16'h0000;
        rom[2][1212] = 16'h0000;
        rom[2][1213] = 16'h0000;
        rom[2][1214] = 16'h0000;
        rom[2][1215] = 16'h0000;
        rom[2][1216] = 16'h0000;
        rom[2][1217] = 16'h0000;
        rom[2][1218] = 16'h0000;
        rom[2][1219] = 16'h0000;
        rom[2][1220] = 16'h0000;
        rom[2][1221] = 16'h0000;
        rom[2][1222] = 16'h0000;
        rom[2][1223] = 16'h0000;
        rom[2][1224] = 16'h0000;
        rom[2][1225] = 16'h0000;
        rom[2][1226] = 16'h0000;
        rom[2][1227] = 16'h0000;
        rom[2][1228] = 16'h0000;
        rom[2][1229] = 16'h0000;
        rom[2][1230] = 16'h0000;
        rom[2][1231] = 16'h0000;
        rom[2][1232] = 16'h0000;
        rom[2][1233] = 16'h0000;
        rom[2][1234] = 16'h0000;
        rom[2][1235] = 16'h0000;
        rom[2][1236] = 16'h0000;
        rom[2][1237] = 16'h0000;
        rom[2][1238] = 16'h0000;
        rom[2][1239] = 16'h0000;
        rom[2][1240] = 16'h0000;
        rom[2][1241] = 16'h0000;
        rom[2][1242] = 16'h0000;
        rom[2][1243] = 16'h0000;
        rom[2][1244] = 16'h0000;
        rom[2][1245] = 16'h0000;
        rom[2][1246] = 16'h0000;
        rom[2][1247] = 16'h0000;
        rom[2][1248] = 16'h0000;
        rom[2][1249] = 16'h0000;
        rom[2][1250] = 16'h0000;
        rom[2][1251] = 16'h0000;
        rom[2][1252] = 16'h0000;
        rom[2][1253] = 16'h0000;
        rom[2][1254] = 16'h0000;
        rom[2][1255] = 16'h0000;
        rom[2][1256] = 16'h0000;
        rom[2][1257] = 16'h0000;
        rom[2][1258] = 16'h0000;
        rom[2][1259] = 16'h0000;
        rom[2][1260] = 16'h0000;
        rom[2][1261] = 16'h0000;
        rom[2][1262] = 16'h0000;
        rom[2][1263] = 16'h0000;
        rom[2][1264] = 16'h0000;
        rom[2][1265] = 16'h0000;
        rom[2][1266] = 16'h0000;
        rom[2][1267] = 16'h0000;
        rom[2][1268] = 16'h0000;
        rom[2][1269] = 16'h0000;
        rom[2][1270] = 16'h0000;
        rom[2][1271] = 16'h0000;
        rom[2][1272] = 16'h0000;
        rom[2][1273] = 16'h0000;
        rom[3][0] = 16'h0121;
        rom[3][1] = 16'h0119;
        rom[3][2] = 16'h0119;
        rom[3][3] = 16'h010B;
        rom[3][4] = 16'h00CA;
        rom[3][5] = 16'h0098;
        rom[3][6] = 16'h0073;
        rom[3][7] = 16'h0048;
        rom[3][8] = 16'h0024;
        rom[3][9] = 16'hFFF9;
        rom[3][10] = 16'hFFE3;
        rom[3][11] = 16'hFFCD;
        rom[3][12] = 16'hFFBF;
        rom[3][13] = 16'hFFA9;
        rom[3][14] = 16'hFF9B;
        rom[3][15] = 16'hFF8D;
        rom[3][16] = 16'hFF8D;
        rom[3][17] = 16'hFF9B;
        rom[3][18] = 16'hFFB8;
        rom[3][19] = 16'h0057;
        rom[3][20] = 16'h00CA;
        rom[3][21] = 16'h00E0;
        rom[3][22] = 16'h010B;
        rom[3][23] = 16'h013E;
        rom[3][24] = 16'h0162;
        rom[3][25] = 16'h0170;
        rom[3][26] = 16'h0136;
        rom[3][27] = 16'h00F5;
        rom[3][28] = 16'h00EE;
        rom[3][29] = 16'h00F5;
        rom[3][30] = 16'h0104;
        rom[3][31] = 16'h00F5;
        rom[3][32] = 16'h0000;
        rom[3][33] = 16'h0000;
        rom[3][34] = 16'h0000;
        rom[3][35] = 16'h0000;
        rom[3][36] = 16'h0000;
        rom[3][37] = 16'h0000;
        rom[3][38] = 16'h0000;
        rom[3][39] = 16'h0000;
        rom[3][40] = 16'h0000;
        rom[3][41] = 16'h0000;
        rom[3][42] = 16'h0000;
        rom[3][43] = 16'h0000;
        rom[3][44] = 16'h0000;
        rom[3][45] = 16'h0000;
        rom[3][46] = 16'h0000;
        rom[3][47] = 16'h0000;
        rom[3][48] = 16'h0000;
        rom[3][49] = 16'h0000;
        rom[3][50] = 16'h0000;
        rom[3][51] = 16'h0000;
        rom[3][52] = 16'h0000;
        rom[3][53] = 16'h0000;
        rom[3][54] = 16'h0000;
        rom[3][55] = 16'h0000;
        rom[3][56] = 16'h0000;
        rom[3][57] = 16'h0000;
        rom[3][58] = 16'h0000;
        rom[3][59] = 16'h0000;
        rom[3][60] = 16'h0000;
        rom[3][61] = 16'h0000;
        rom[3][62] = 16'h0000;
        rom[3][63] = 16'h0000;
        rom[3][64] = 16'h0000;
        rom[3][65] = 16'h0000;
        rom[3][66] = 16'h0000;
        rom[3][67] = 16'h0000;
        rom[3][68] = 16'h0000;
        rom[3][69] = 16'h0000;
        rom[3][70] = 16'h0000;
        rom[3][71] = 16'h0000;
        rom[3][72] = 16'h0000;
        rom[3][73] = 16'h0000;
        rom[3][74] = 16'h0000;
        rom[3][75] = 16'h0000;
        rom[3][76] = 16'h0000;
        rom[3][77] = 16'h0000;
        rom[3][78] = 16'h0000;
        rom[3][79] = 16'h0000;
        rom[3][80] = 16'h0000;
        rom[3][81] = 16'h0000;
        rom[3][82] = 16'h0000;
        rom[3][83] = 16'h0000;
        rom[3][84] = 16'h0000;
        rom[3][85] = 16'h0000;
        rom[3][86] = 16'h0000;
        rom[3][87] = 16'h0000;
        rom[3][88] = 16'h0000;
        rom[3][89] = 16'h0000;
        rom[3][90] = 16'h0000;
        rom[3][91] = 16'h0000;
        rom[3][92] = 16'h0000;
        rom[3][93] = 16'h0000;
        rom[3][94] = 16'h0000;
        rom[3][95] = 16'h0000;
        rom[3][96] = 16'h0000;
        rom[3][97] = 16'h0000;
        rom[3][98] = 16'h001D;
        rom[3][99] = 16'h000E;
        rom[3][100] = 16'hFFBF;
        rom[3][101] = 16'hFF7E;
        rom[3][102] = 16'hFF9B;
        rom[3][103] = 16'hFFB1;
        rom[3][104] = 16'hFF8D;
        rom[3][105] = 16'hFF5A;
        rom[3][106] = 16'hFF36;
        rom[3][107] = 16'hFF61;
        rom[3][108] = 16'hFF53;
        rom[3][109] = 16'hFF44;
        rom[3][110] = 16'hFF44;
        rom[3][111] = 16'hFF2F;
        rom[3][112] = 16'hFF2F;
        rom[3][113] = 16'hFF20;
        rom[3][114] = 16'hFF2F;
        rom[3][115] = 16'hFF53;
        rom[3][116] = 16'hFF7E;
        rom[3][117] = 16'hFF85;
        rom[3][118] = 16'hFF68;
        rom[3][119] = 16'hFF53;
        rom[3][120] = 16'hFF8D;
        rom[3][121] = 16'hFFEA;
        rom[3][122] = 16'h0033;
        rom[3][123] = 16'h0065;
        rom[3][124] = 16'h006C;
        rom[3][125] = 16'h005E;
        rom[3][126] = 16'h0048;
        rom[3][127] = 16'h003A;
        rom[3][128] = 16'h000E;
        rom[3][129] = 16'hFFF9;
        rom[3][130] = 16'h0000;
        rom[3][131] = 16'h0000;
        rom[3][132] = 16'h0000;
        rom[3][133] = 16'h0000;
        rom[3][134] = 16'h0000;
        rom[3][135] = 16'h0000;
        rom[3][136] = 16'h0000;
        rom[3][137] = 16'h0000;
        rom[3][138] = 16'h0000;
        rom[3][139] = 16'h0000;
        rom[3][140] = 16'h0000;
        rom[3][141] = 16'h0000;
        rom[3][142] = 16'h0000;
        rom[3][143] = 16'h0000;
        rom[3][144] = 16'h0000;
        rom[3][145] = 16'h0000;
        rom[3][146] = 16'h0000;
        rom[3][147] = 16'h0000;
        rom[3][148] = 16'h0000;
        rom[3][149] = 16'h0000;
        rom[3][150] = 16'h0000;
        rom[3][151] = 16'h0000;
        rom[3][152] = 16'h0000;
        rom[3][153] = 16'h0000;
        rom[3][154] = 16'h0000;
        rom[3][155] = 16'h0000;
        rom[3][156] = 16'h0000;
        rom[3][157] = 16'h0000;
        rom[3][158] = 16'h0000;
        rom[3][159] = 16'h0000;
        rom[3][160] = 16'h0000;
        rom[3][161] = 16'h0000;
        rom[3][162] = 16'h0000;
        rom[3][163] = 16'h0000;
        rom[3][164] = 16'h0000;
        rom[3][165] = 16'h0000;
        rom[3][166] = 16'h0000;
        rom[3][167] = 16'h0000;
        rom[3][168] = 16'h0000;
        rom[3][169] = 16'h0000;
        rom[3][170] = 16'h0000;
        rom[3][171] = 16'h0000;
        rom[3][172] = 16'h0000;
        rom[3][173] = 16'h0000;
        rom[3][174] = 16'h0000;
        rom[3][175] = 16'h0000;
        rom[3][176] = 16'h0000;
        rom[3][177] = 16'h0000;
        rom[3][178] = 16'h0000;
        rom[3][179] = 16'h0000;
        rom[3][180] = 16'h0000;
        rom[3][181] = 16'h0000;
        rom[3][182] = 16'h0000;
        rom[3][183] = 16'h0000;
        rom[3][184] = 16'h0000;
        rom[3][185] = 16'h0000;
        rom[3][186] = 16'h0000;
        rom[3][187] = 16'h0000;
        rom[3][188] = 16'h0000;
        rom[3][189] = 16'h0000;
        rom[3][190] = 16'h0000;
        rom[3][191] = 16'h0000;
        rom[3][192] = 16'h0000;
        rom[3][193] = 16'h0000;
        rom[3][194] = 16'h0000;
        rom[3][195] = 16'h0000;
        rom[3][196] = 16'hFFEA;
        rom[3][197] = 16'h0007;
        rom[3][198] = 16'h0007;
        rom[3][199] = 16'h001D;
        rom[3][200] = 16'h0000;
        rom[3][201] = 16'hFFF2;
        rom[3][202] = 16'h0000;
        rom[3][203] = 16'h007B;
        rom[3][204] = 16'h0082;
        rom[3][205] = 16'h003A;
        rom[3][206] = 16'h0041;
        rom[3][207] = 16'h004F;
        rom[3][208] = 16'h0041;
        rom[3][209] = 16'h0048;
        rom[3][210] = 16'h0033;
        rom[3][211] = 16'h0033;
        rom[3][212] = 16'h0057;
        rom[3][213] = 16'h0089;
        rom[3][214] = 16'h00A6;
        rom[3][215] = 16'h000E;
        rom[3][216] = 16'hFFA9;
        rom[3][217] = 16'hFF68;
        rom[3][218] = 16'hFED1;
        rom[3][219] = 16'hFE56;
        rom[3][220] = 16'hFE39;
        rom[3][221] = 16'hFE89;
        rom[3][222] = 16'hFF4C;
        rom[3][223] = 16'h004F;
        rom[3][224] = 16'h0090;
        rom[3][225] = 16'h0082;
        rom[3][226] = 16'h0033;
        rom[3][227] = 16'hFFEA;
        rom[3][228] = 16'h0000;
        rom[3][229] = 16'h0000;
        rom[3][230] = 16'h0000;
        rom[3][231] = 16'h0000;
        rom[3][232] = 16'h0000;
        rom[3][233] = 16'h0000;
        rom[3][234] = 16'h0000;
        rom[3][235] = 16'h0000;
        rom[3][236] = 16'h0000;
        rom[3][237] = 16'h0000;
        rom[3][238] = 16'h0000;
        rom[3][239] = 16'h0000;
        rom[3][240] = 16'h0000;
        rom[3][241] = 16'h0000;
        rom[3][242] = 16'h0000;
        rom[3][243] = 16'h0000;
        rom[3][244] = 16'h0000;
        rom[3][245] = 16'h0000;
        rom[3][246] = 16'h0000;
        rom[3][247] = 16'h0000;
        rom[3][248] = 16'h0000;
        rom[3][249] = 16'h0000;
        rom[3][250] = 16'h0000;
        rom[3][251] = 16'h0000;
        rom[3][252] = 16'h0000;
        rom[3][253] = 16'h0000;
        rom[3][254] = 16'h0000;
        rom[3][255] = 16'h0000;
        rom[3][256] = 16'h0000;
        rom[3][257] = 16'h0000;
        rom[3][258] = 16'h0000;
        rom[3][259] = 16'h0000;
        rom[3][260] = 16'h0000;
        rom[3][261] = 16'h0000;
        rom[3][262] = 16'h0000;
        rom[3][263] = 16'h0000;
        rom[3][264] = 16'h0000;
        rom[3][265] = 16'h0000;
        rom[3][266] = 16'h0000;
        rom[3][267] = 16'h0000;
        rom[3][268] = 16'h0000;
        rom[3][269] = 16'h0000;
        rom[3][270] = 16'h0000;
        rom[3][271] = 16'h0000;
        rom[3][272] = 16'h0000;
        rom[3][273] = 16'h0000;
        rom[3][274] = 16'h0000;
        rom[3][275] = 16'h0000;
        rom[3][276] = 16'h0000;
        rom[3][277] = 16'h0000;
        rom[3][278] = 16'h0000;
        rom[3][279] = 16'h0000;
        rom[3][280] = 16'h0000;
        rom[3][281] = 16'h0000;
        rom[3][282] = 16'h0000;
        rom[3][283] = 16'h0000;
        rom[3][284] = 16'h0000;
        rom[3][285] = 16'h0000;
        rom[3][286] = 16'h0000;
        rom[3][287] = 16'h0000;
        rom[3][288] = 16'h0000;
        rom[3][289] = 16'h0000;
        rom[3][290] = 16'h0000;
        rom[3][291] = 16'h0000;
        rom[3][292] = 16'h0000;
        rom[3][293] = 16'h0000;
        rom[3][294] = 16'h0082;
        rom[3][295] = 16'h0082;
        rom[3][296] = 16'h00C3;
        rom[3][297] = 16'h00C3;
        rom[3][298] = 16'h0082;
        rom[3][299] = 16'h0089;
        rom[3][300] = 16'h0073;
        rom[3][301] = 16'hFFF9;
        rom[3][302] = 16'hFFDC;
        rom[3][303] = 16'h0007;
        rom[3][304] = 16'h000E;
        rom[3][305] = 16'h0016;
        rom[3][306] = 16'h0024;
        rom[3][307] = 16'h0041;
        rom[3][308] = 16'h0033;
        rom[3][309] = 16'h0024;
        rom[3][310] = 16'h0048;
        rom[3][311] = 16'h007B;
        rom[3][312] = 16'h00B4;
        rom[3][313] = 16'h0121;
        rom[3][314] = 16'h0162;
        rom[3][315] = 16'h0121;
        rom[3][316] = 16'h00D1;
        rom[3][317] = 16'h0024;
        rom[3][318] = 16'hFFD5;
        rom[3][319] = 16'hFFA2;
        rom[3][320] = 16'hFF77;
        rom[3][321] = 16'hFFEA;
        rom[3][322] = 16'h0089;
        rom[3][323] = 16'h00D9;
        rom[3][324] = 16'h00E7;
        rom[3][325] = 16'h00B4;
        rom[3][326] = 16'h0000;
        rom[3][327] = 16'h0000;
        rom[3][328] = 16'h0000;
        rom[3][329] = 16'h0000;
        rom[3][330] = 16'h0000;
        rom[3][331] = 16'h0000;
        rom[3][332] = 16'h0000;
        rom[3][333] = 16'h0000;
        rom[3][334] = 16'h0000;
        rom[3][335] = 16'h0000;
        rom[3][336] = 16'h0000;
        rom[3][337] = 16'h0000;
        rom[3][338] = 16'h0000;
        rom[3][339] = 16'h0000;
        rom[3][340] = 16'h0000;
        rom[3][341] = 16'h0000;
        rom[3][342] = 16'h0000;
        rom[3][343] = 16'h0000;
        rom[3][344] = 16'h0000;
        rom[3][345] = 16'h0000;
        rom[3][346] = 16'h0000;
        rom[3][347] = 16'h0000;
        rom[3][348] = 16'h0000;
        rom[3][349] = 16'h0000;
        rom[3][350] = 16'h0000;
        rom[3][351] = 16'h0000;
        rom[3][352] = 16'h0000;
        rom[3][353] = 16'h0000;
        rom[3][354] = 16'h0000;
        rom[3][355] = 16'h0000;
        rom[3][356] = 16'h0000;
        rom[3][357] = 16'h0000;
        rom[3][358] = 16'h0000;
        rom[3][359] = 16'h0000;
        rom[3][360] = 16'h0000;
        rom[3][361] = 16'h0000;
        rom[3][362] = 16'h0000;
        rom[3][363] = 16'h0000;
        rom[3][364] = 16'h0000;
        rom[3][365] = 16'h0000;
        rom[3][366] = 16'h0000;
        rom[3][367] = 16'h0000;
        rom[3][368] = 16'h0000;
        rom[3][369] = 16'h0000;
        rom[3][370] = 16'h0000;
        rom[3][371] = 16'h0000;
        rom[3][372] = 16'h0000;
        rom[3][373] = 16'h0000;
        rom[3][374] = 16'h0000;
        rom[3][375] = 16'h0000;
        rom[3][376] = 16'h0000;
        rom[3][377] = 16'h0000;
        rom[3][378] = 16'h0000;
        rom[3][379] = 16'h0000;
        rom[3][380] = 16'h0000;
        rom[3][381] = 16'h0000;
        rom[3][382] = 16'h0000;
        rom[3][383] = 16'h0000;
        rom[3][384] = 16'h0000;
        rom[3][385] = 16'h0000;
        rom[3][386] = 16'h0000;
        rom[3][387] = 16'h0000;
        rom[3][388] = 16'h0000;
        rom[3][389] = 16'h0000;
        rom[3][390] = 16'h0000;
        rom[3][391] = 16'h0000;
        rom[3][392] = 16'h001D;
        rom[3][393] = 16'hFFF2;
        rom[3][394] = 16'hFFB1;
        rom[3][395] = 16'hFFBF;
        rom[3][396] = 16'h000E;
        rom[3][397] = 16'h000E;
        rom[3][398] = 16'h001D;
        rom[3][399] = 16'h0065;
        rom[3][400] = 16'h0057;
        rom[3][401] = 16'h003A;
        rom[3][402] = 16'h003A;
        rom[3][403] = 16'h0065;
        rom[3][404] = 16'h0090;
        rom[3][405] = 16'h00AD;
        rom[3][406] = 16'h0090;
        rom[3][407] = 16'h0089;
        rom[3][408] = 16'h00AD;
        rom[3][409] = 16'h00C3;
        rom[3][410] = 16'h00B4;
        rom[3][411] = 16'hFFEA;
        rom[3][412] = 16'hFF53;
        rom[3][413] = 16'hFF20;
        rom[3][414] = 16'hFF77;
        rom[3][415] = 16'hFF77;
        rom[3][416] = 16'hFF2F;
        rom[3][417] = 16'hFED8;
        rom[3][418] = 16'hFE73;
        rom[3][419] = 16'hFEBB;
        rom[3][420] = 16'hFF3D;
        rom[3][421] = 16'hFF7E;
        rom[3][422] = 16'hFFE3;
        rom[3][423] = 16'hFF7E;
        rom[3][424] = 16'h0000;
        rom[3][425] = 16'h0000;
        rom[3][426] = 16'h0000;
        rom[3][427] = 16'h0000;
        rom[3][428] = 16'h0000;
        rom[3][429] = 16'h0000;
        rom[3][430] = 16'h0000;
        rom[3][431] = 16'h0000;
        rom[3][432] = 16'h0000;
        rom[3][433] = 16'h0000;
        rom[3][434] = 16'h0000;
        rom[3][435] = 16'h0000;
        rom[3][436] = 16'h0000;
        rom[3][437] = 16'h0000;
        rom[3][438] = 16'h0000;
        rom[3][439] = 16'h0000;
        rom[3][440] = 16'h0000;
        rom[3][441] = 16'h0000;
        rom[3][442] = 16'h0000;
        rom[3][443] = 16'h0000;
        rom[3][444] = 16'h0000;
        rom[3][445] = 16'h0000;
        rom[3][446] = 16'h0000;
        rom[3][447] = 16'h0000;
        rom[3][448] = 16'h0000;
        rom[3][449] = 16'h0000;
        rom[3][450] = 16'h0000;
        rom[3][451] = 16'h0000;
        rom[3][452] = 16'h0000;
        rom[3][453] = 16'h0000;
        rom[3][454] = 16'h0000;
        rom[3][455] = 16'h0000;
        rom[3][456] = 16'h0000;
        rom[3][457] = 16'h0000;
        rom[3][458] = 16'h0000;
        rom[3][459] = 16'h0000;
        rom[3][460] = 16'h0000;
        rom[3][461] = 16'h0000;
        rom[3][462] = 16'h0000;
        rom[3][463] = 16'h0000;
        rom[3][464] = 16'h0000;
        rom[3][465] = 16'h0000;
        rom[3][466] = 16'h0000;
        rom[3][467] = 16'h0000;
        rom[3][468] = 16'h0000;
        rom[3][469] = 16'h0000;
        rom[3][470] = 16'h0000;
        rom[3][471] = 16'h0000;
        rom[3][472] = 16'h0000;
        rom[3][473] = 16'h0000;
        rom[3][474] = 16'h0000;
        rom[3][475] = 16'h0000;
        rom[3][476] = 16'h0000;
        rom[3][477] = 16'h0000;
        rom[3][478] = 16'h0000;
        rom[3][479] = 16'h0000;
        rom[3][480] = 16'h0000;
        rom[3][481] = 16'h0000;
        rom[3][482] = 16'h0000;
        rom[3][483] = 16'h0000;
        rom[3][484] = 16'h0000;
        rom[3][485] = 16'h0000;
        rom[3][486] = 16'h0000;
        rom[3][487] = 16'h0000;
        rom[3][488] = 16'h0000;
        rom[3][489] = 16'h0000;
        rom[3][490] = 16'h000E;
        rom[3][491] = 16'hFFF2;
        rom[3][492] = 16'h0073;
        rom[3][493] = 16'h009F;
        rom[3][494] = 16'h00A6;
        rom[3][495] = 16'h00CA;
        rom[3][496] = 16'h00D9;
        rom[3][497] = 16'h0090;
        rom[3][498] = 16'h006C;
        rom[3][499] = 16'h00A6;
        rom[3][500] = 16'h00B4;
        rom[3][501] = 16'h0082;
        rom[3][502] = 16'h009F;
        rom[3][503] = 16'h00E0;
        rom[3][504] = 16'h00E7;
        rom[3][505] = 16'h00CA;
        rom[3][506] = 16'h00E0;
        rom[3][507] = 16'h00D9;
        rom[3][508] = 16'h0065;
        rom[3][509] = 16'h0048;
        rom[3][510] = 16'h0065;
        rom[3][511] = 16'h0089;
        rom[3][512] = 16'h0090;
        rom[3][513] = 16'h0082;
        rom[3][514] = 16'h00EE;
        rom[3][515] = 16'h014C;
        rom[3][516] = 16'h0153;
        rom[3][517] = 16'h005E;
        rom[3][518] = 16'hFFD5;
        rom[3][519] = 16'hFFF2;
        rom[3][520] = 16'h0089;
        rom[3][521] = 16'h006C;
        rom[3][522] = 16'h0000;
        rom[3][523] = 16'h0000;
        rom[3][524] = 16'h0000;
        rom[3][525] = 16'h0000;
        rom[3][526] = 16'h0000;
        rom[3][527] = 16'h0000;
        rom[3][528] = 16'h0000;
        rom[3][529] = 16'h0000;
        rom[3][530] = 16'h0000;
        rom[3][531] = 16'h0000;
        rom[3][532] = 16'h0000;
        rom[3][533] = 16'h0000;
        rom[3][534] = 16'h0000;
        rom[3][535] = 16'h0000;
        rom[3][536] = 16'h0000;
        rom[3][537] = 16'h0000;
        rom[3][538] = 16'h0000;
        rom[3][539] = 16'h0000;
        rom[3][540] = 16'h0000;
        rom[3][541] = 16'h0000;
        rom[3][542] = 16'h0000;
        rom[3][543] = 16'h0000;
        rom[3][544] = 16'h0000;
        rom[3][545] = 16'h0000;
        rom[3][546] = 16'h0000;
        rom[3][547] = 16'h0000;
        rom[3][548] = 16'h0000;
        rom[3][549] = 16'h0000;
        rom[3][550] = 16'h0000;
        rom[3][551] = 16'h0000;
        rom[3][552] = 16'h0000;
        rom[3][553] = 16'h0000;
        rom[3][554] = 16'h0000;
        rom[3][555] = 16'h0000;
        rom[3][556] = 16'h0000;
        rom[3][557] = 16'h0000;
        rom[3][558] = 16'h0000;
        rom[3][559] = 16'h0000;
        rom[3][560] = 16'h0000;
        rom[3][561] = 16'h0000;
        rom[3][562] = 16'h0000;
        rom[3][563] = 16'h0000;
        rom[3][564] = 16'h0000;
        rom[3][565] = 16'h0000;
        rom[3][566] = 16'h0000;
        rom[3][567] = 16'h0000;
        rom[3][568] = 16'h0000;
        rom[3][569] = 16'h0000;
        rom[3][570] = 16'h0000;
        rom[3][571] = 16'h0000;
        rom[3][572] = 16'h0000;
        rom[3][573] = 16'h0000;
        rom[3][574] = 16'h0000;
        rom[3][575] = 16'h0000;
        rom[3][576] = 16'h0000;
        rom[3][577] = 16'h0000;
        rom[3][578] = 16'h0000;
        rom[3][579] = 16'h0000;
        rom[3][580] = 16'h0000;
        rom[3][581] = 16'h0000;
        rom[3][582] = 16'h0000;
        rom[3][583] = 16'h0000;
        rom[3][584] = 16'h0000;
        rom[3][585] = 16'h0000;
        rom[3][586] = 16'h0000;
        rom[3][587] = 16'h0000;
        rom[3][588] = 16'hFFEA;
        rom[3][589] = 16'hFFD5;
        rom[3][590] = 16'hFF70;
        rom[3][591] = 16'hFFC6;
        rom[3][592] = 16'h0016;
        rom[3][593] = 16'h0033;
        rom[3][594] = 16'hFFF2;
        rom[3][595] = 16'h000E;
        rom[3][596] = 16'hFFF9;
        rom[3][597] = 16'h0016;
        rom[3][598] = 16'h0016;
        rom[3][599] = 16'hFFEA;
        rom[3][600] = 16'h0048;
        rom[3][601] = 16'h004F;
        rom[3][602] = 16'h005E;
        rom[3][603] = 16'h0065;
        rom[3][604] = 16'h003A;
        rom[3][605] = 16'h0073;
        rom[3][606] = 16'h0033;
        rom[3][607] = 16'hFF44;
        rom[3][608] = 16'hFED1;
        rom[3][609] = 16'hFEE7;
        rom[3][610] = 16'hFED1;
        rom[3][611] = 16'hFEAD;
        rom[3][612] = 16'hFED1;
        rom[3][613] = 16'hFF7E;
        rom[3][614] = 16'h005E;
        rom[3][615] = 16'h0024;
        rom[3][616] = 16'hFFA2;
        rom[3][617] = 16'hFF9B;
        rom[3][618] = 16'hFFE3;
        rom[3][619] = 16'h0024;
        rom[3][620] = 16'h0000;
        rom[3][621] = 16'h0000;
        rom[3][622] = 16'h0000;
        rom[3][623] = 16'h0000;
        rom[3][624] = 16'h0000;
        rom[3][625] = 16'h0000;
        rom[3][626] = 16'h0000;
        rom[3][627] = 16'h0000;
        rom[3][628] = 16'h0000;
        rom[3][629] = 16'h0000;
        rom[3][630] = 16'h0000;
        rom[3][631] = 16'h0000;
        rom[3][632] = 16'h0000;
        rom[3][633] = 16'h0000;
        rom[3][634] = 16'h0000;
        rom[3][635] = 16'h0000;
        rom[3][636] = 16'h0000;
        rom[3][637] = 16'h0000;
        rom[3][638] = 16'h0000;
        rom[3][639] = 16'h0000;
        rom[3][640] = 16'h0000;
        rom[3][641] = 16'h0000;
        rom[3][642] = 16'h0000;
        rom[3][643] = 16'h0000;
        rom[3][644] = 16'h0000;
        rom[3][645] = 16'h0000;
        rom[3][646] = 16'h0000;
        rom[3][647] = 16'h0000;
        rom[3][648] = 16'h0000;
        rom[3][649] = 16'h0000;
        rom[3][650] = 16'h0000;
        rom[3][651] = 16'h0000;
        rom[3][652] = 16'h0000;
        rom[3][653] = 16'h0000;
        rom[3][654] = 16'h0000;
        rom[3][655] = 16'h0000;
        rom[3][656] = 16'h0000;
        rom[3][657] = 16'h0000;
        rom[3][658] = 16'h0000;
        rom[3][659] = 16'h0000;
        rom[3][660] = 16'h0000;
        rom[3][661] = 16'h0000;
        rom[3][662] = 16'h0000;
        rom[3][663] = 16'h0000;
        rom[3][664] = 16'h0000;
        rom[3][665] = 16'h0000;
        rom[3][666] = 16'h0000;
        rom[3][667] = 16'h0000;
        rom[3][668] = 16'h0000;
        rom[3][669] = 16'h0000;
        rom[3][670] = 16'h0000;
        rom[3][671] = 16'h0000;
        rom[3][672] = 16'h0000;
        rom[3][673] = 16'h0000;
        rom[3][674] = 16'h0000;
        rom[3][675] = 16'h0000;
        rom[3][676] = 16'h0000;
        rom[3][677] = 16'h0000;
        rom[3][678] = 16'h0000;
        rom[3][679] = 16'h0000;
        rom[3][680] = 16'h0000;
        rom[3][681] = 16'h0000;
        rom[3][682] = 16'h0000;
        rom[3][683] = 16'h0000;
        rom[3][684] = 16'h0000;
        rom[3][685] = 16'h0000;
        rom[3][686] = 16'h0119;
        rom[3][687] = 16'h00D1;
        rom[3][688] = 16'h00FD;
        rom[3][689] = 16'h010B;
        rom[3][690] = 16'h00FD;
        rom[3][691] = 16'h00D9;
        rom[3][692] = 16'h0082;
        rom[3][693] = 16'h009F;
        rom[3][694] = 16'h00D9;
        rom[3][695] = 16'h00F5;
        rom[3][696] = 16'h00D1;
        rom[3][697] = 16'h00E0;
        rom[3][698] = 16'h00F5;
        rom[3][699] = 16'h00A6;
        rom[3][700] = 16'h00A6;
        rom[3][701] = 16'h00D1;
        rom[3][702] = 16'h00C3;
        rom[3][703] = 16'h00D1;
        rom[3][704] = 16'h00C3;
        rom[3][705] = 16'h00B4;
        rom[3][706] = 16'h00D1;
        rom[3][707] = 16'h00BC;
        rom[3][708] = 16'h0082;
        rom[3][709] = 16'hFFCD;
        rom[3][710] = 16'hFEEE;
        rom[3][711] = 16'hFEAD;
        rom[3][712] = 16'hFF44;
        rom[3][713] = 16'h009F;
        rom[3][714] = 16'h00C3;
        rom[3][715] = 16'h00BC;
        rom[3][716] = 16'h009F;
        rom[3][717] = 16'h00E7;
        rom[3][718] = 16'h0000;
        rom[3][719] = 16'h0000;
        rom[3][720] = 16'h0000;
        rom[3][721] = 16'h0000;
        rom[3][722] = 16'h0000;
        rom[3][723] = 16'h0000;
        rom[3][724] = 16'h0000;
        rom[3][725] = 16'h0000;
        rom[3][726] = 16'h0000;
        rom[3][727] = 16'h0000;
        rom[3][728] = 16'h0000;
        rom[3][729] = 16'h0000;
        rom[3][730] = 16'h0000;
        rom[3][731] = 16'h0000;
        rom[3][732] = 16'h0000;
        rom[3][733] = 16'h0000;
        rom[3][734] = 16'h0000;
        rom[3][735] = 16'h0000;
        rom[3][736] = 16'h0000;
        rom[3][737] = 16'h0000;
        rom[3][738] = 16'h0000;
        rom[3][739] = 16'h0000;
        rom[3][740] = 16'h0000;
        rom[3][741] = 16'h0000;
        rom[3][742] = 16'h0000;
        rom[3][743] = 16'h0000;
        rom[3][744] = 16'h0000;
        rom[3][745] = 16'h0000;
        rom[3][746] = 16'h0000;
        rom[3][747] = 16'h0000;
        rom[3][748] = 16'h0000;
        rom[3][749] = 16'h0000;
        rom[3][750] = 16'h0000;
        rom[3][751] = 16'h0000;
        rom[3][752] = 16'h0000;
        rom[3][753] = 16'h0000;
        rom[3][754] = 16'h0000;
        rom[3][755] = 16'h0000;
        rom[3][756] = 16'h0000;
        rom[3][757] = 16'h0000;
        rom[3][758] = 16'h0000;
        rom[3][759] = 16'h0000;
        rom[3][760] = 16'h0000;
        rom[3][761] = 16'h0000;
        rom[3][762] = 16'h0000;
        rom[3][763] = 16'h0000;
        rom[3][764] = 16'h0000;
        rom[3][765] = 16'h0000;
        rom[3][766] = 16'h0000;
        rom[3][767] = 16'h0000;
        rom[3][768] = 16'h0000;
        rom[3][769] = 16'h0000;
        rom[3][770] = 16'h0000;
        rom[3][771] = 16'h0000;
        rom[3][772] = 16'h0000;
        rom[3][773] = 16'h0000;
        rom[3][774] = 16'h0000;
        rom[3][775] = 16'h0000;
        rom[3][776] = 16'h0000;
        rom[3][777] = 16'h0000;
        rom[3][778] = 16'h0000;
        rom[3][779] = 16'h0000;
        rom[3][780] = 16'h0000;
        rom[3][781] = 16'h0000;
        rom[3][782] = 16'h0000;
        rom[3][783] = 16'h0000;
        rom[3][784] = 16'h005E;
        rom[3][785] = 16'hFFEA;
        rom[3][786] = 16'hFFDC;
        rom[3][787] = 16'h0048;
        rom[3][788] = 16'h003A;
        rom[3][789] = 16'h0041;
        rom[3][790] = 16'h003A;
        rom[3][791] = 16'hFF7E;
        rom[3][792] = 16'hFFF9;
        rom[3][793] = 16'h0089;
        rom[3][794] = 16'h0065;
        rom[3][795] = 16'h005E;
        rom[3][796] = 16'h0057;
        rom[3][797] = 16'h0048;
        rom[3][798] = 16'h007B;
        rom[3][799] = 16'h0057;
        rom[3][800] = 16'h0033;
        rom[3][801] = 16'h005E;
        rom[3][802] = 16'h000E;
        rom[3][803] = 16'h004F;
        rom[3][804] = 16'h006C;
        rom[3][805] = 16'h009F;
        rom[3][806] = 16'h014C;
        rom[3][807] = 16'h00EE;
        rom[3][808] = 16'h004F;
        rom[3][809] = 16'hFF94;
        rom[3][810] = 16'hFF3D;
        rom[3][811] = 16'hFFDC;
        rom[3][812] = 16'h003A;
        rom[3][813] = 16'hFFEA;
        rom[3][814] = 16'hFF53;
        rom[3][815] = 16'hFF36;
        rom[3][816] = 16'h0000;
        rom[3][817] = 16'h0000;
        rom[3][818] = 16'h0000;
        rom[3][819] = 16'h0000;
        rom[3][820] = 16'h0000;
        rom[3][821] = 16'h0000;
        rom[3][822] = 16'h0000;
        rom[3][823] = 16'h0000;
        rom[3][824] = 16'h0000;
        rom[3][825] = 16'h0000;
        rom[3][826] = 16'h0000;
        rom[3][827] = 16'h0000;
        rom[3][828] = 16'h0000;
        rom[3][829] = 16'h0000;
        rom[3][830] = 16'h0000;
        rom[3][831] = 16'h0000;
        rom[3][832] = 16'h0000;
        rom[3][833] = 16'h0000;
        rom[3][834] = 16'h0000;
        rom[3][835] = 16'h0000;
        rom[3][836] = 16'h0000;
        rom[3][837] = 16'h0000;
        rom[3][838] = 16'h0000;
        rom[3][839] = 16'h0000;
        rom[3][840] = 16'h0000;
        rom[3][841] = 16'h0000;
        rom[3][842] = 16'h0000;
        rom[3][843] = 16'h0000;
        rom[3][844] = 16'h0000;
        rom[3][845] = 16'h0000;
        rom[3][846] = 16'h0000;
        rom[3][847] = 16'h0000;
        rom[3][848] = 16'h0000;
        rom[3][849] = 16'h0000;
        rom[3][850] = 16'h0000;
        rom[3][851] = 16'h0000;
        rom[3][852] = 16'h0000;
        rom[3][853] = 16'h0000;
        rom[3][854] = 16'h0000;
        rom[3][855] = 16'h0000;
        rom[3][856] = 16'h0000;
        rom[3][857] = 16'h0000;
        rom[3][858] = 16'h0000;
        rom[3][859] = 16'h0000;
        rom[3][860] = 16'h0000;
        rom[3][861] = 16'h0000;
        rom[3][862] = 16'h0000;
        rom[3][863] = 16'h0000;
        rom[3][864] = 16'h0000;
        rom[3][865] = 16'h0000;
        rom[3][866] = 16'h0000;
        rom[3][867] = 16'h0000;
        rom[3][868] = 16'h0000;
        rom[3][869] = 16'h0000;
        rom[3][870] = 16'h0000;
        rom[3][871] = 16'h0000;
        rom[3][872] = 16'h0000;
        rom[3][873] = 16'h0000;
        rom[3][874] = 16'h0000;
        rom[3][875] = 16'h0000;
        rom[3][876] = 16'h0000;
        rom[3][877] = 16'h0000;
        rom[3][878] = 16'h0000;
        rom[3][879] = 16'h0000;
        rom[3][880] = 16'h0000;
        rom[3][881] = 16'h0000;
        rom[3][882] = 16'h0177;
        rom[3][883] = 16'h0112;
        rom[3][884] = 16'h0007;
        rom[3][885] = 16'hFFBF;
        rom[3][886] = 16'h00BC;
        rom[3][887] = 16'h00BC;
        rom[3][888] = 16'h0048;
        rom[3][889] = 16'h0089;
        rom[3][890] = 16'h0104;
        rom[3][891] = 16'h00E0;
        rom[3][892] = 16'h00F5;
        rom[3][893] = 16'h00BC;
        rom[3][894] = 16'h00D9;
        rom[3][895] = 16'h00EE;
        rom[3][896] = 16'h0104;
        rom[3][897] = 16'h00E7;
        rom[3][898] = 16'h00C3;
        rom[3][899] = 16'h009F;
        rom[3][900] = 16'h001D;
        rom[3][901] = 16'hFFDC;
        rom[3][902] = 16'h003A;
        rom[3][903] = 16'h006C;
        rom[3][904] = 16'h0119;
        rom[3][905] = 16'h0186;
        rom[3][906] = 16'h0186;
        rom[3][907] = 16'h015A;
        rom[3][908] = 16'h0089;
        rom[3][909] = 16'h0024;
        rom[3][910] = 16'h00E0;
        rom[3][911] = 16'h015A;
        rom[3][912] = 16'h0104;
        rom[3][913] = 16'h00E0;
        rom[3][914] = 16'h0000;
        rom[3][915] = 16'h0000;
        rom[3][916] = 16'h0000;
        rom[3][917] = 16'h0000;
        rom[3][918] = 16'h0000;
        rom[3][919] = 16'h0000;
        rom[3][920] = 16'h0000;
        rom[3][921] = 16'h0000;
        rom[3][922] = 16'h0000;
        rom[3][923] = 16'h0000;
        rom[3][924] = 16'h0000;
        rom[3][925] = 16'h0000;
        rom[3][926] = 16'h0000;
        rom[3][927] = 16'h0000;
        rom[3][928] = 16'h0000;
        rom[3][929] = 16'h0000;
        rom[3][930] = 16'h0000;
        rom[3][931] = 16'h0000;
        rom[3][932] = 16'h0000;
        rom[3][933] = 16'h0000;
        rom[3][934] = 16'h0000;
        rom[3][935] = 16'h0000;
        rom[3][936] = 16'h0000;
        rom[3][937] = 16'h0000;
        rom[3][938] = 16'h0000;
        rom[3][939] = 16'h0000;
        rom[3][940] = 16'h0000;
        rom[3][941] = 16'h0000;
        rom[3][942] = 16'h0000;
        rom[3][943] = 16'h0000;
        rom[3][944] = 16'h0000;
        rom[3][945] = 16'h0000;
        rom[3][946] = 16'h0000;
        rom[3][947] = 16'h0000;
        rom[3][948] = 16'h0000;
        rom[3][949] = 16'h0000;
        rom[3][950] = 16'h0000;
        rom[3][951] = 16'h0000;
        rom[3][952] = 16'h0000;
        rom[3][953] = 16'h0000;
        rom[3][954] = 16'h0000;
        rom[3][955] = 16'h0000;
        rom[3][956] = 16'h0000;
        rom[3][957] = 16'h0000;
        rom[3][958] = 16'h0000;
        rom[3][959] = 16'h0000;
        rom[3][960] = 16'h0000;
        rom[3][961] = 16'h0000;
        rom[3][962] = 16'h0000;
        rom[3][963] = 16'h0000;
        rom[3][964] = 16'h0000;
        rom[3][965] = 16'h0000;
        rom[3][966] = 16'h0000;
        rom[3][967] = 16'h0000;
        rom[3][968] = 16'h0000;
        rom[3][969] = 16'h0000;
        rom[3][970] = 16'h0000;
        rom[3][971] = 16'h0000;
        rom[3][972] = 16'h0000;
        rom[3][973] = 16'h0000;
        rom[3][974] = 16'h0000;
        rom[3][975] = 16'h0000;
        rom[3][976] = 16'h0000;
        rom[3][977] = 16'h0000;
        rom[3][978] = 16'h0000;
        rom[3][979] = 16'h0000;
        rom[3][980] = 16'h00A6;
        rom[3][981] = 16'h0048;
        rom[3][982] = 16'h0090;
        rom[3][983] = 16'h0112;
        rom[3][984] = 16'h0090;
        rom[3][985] = 16'h000E;
        rom[3][986] = 16'hFFCD;
        rom[3][987] = 16'hFF9B;
        rom[3][988] = 16'hFFF2;
        rom[3][989] = 16'h002B;
        rom[3][990] = 16'h0007;
        rom[3][991] = 16'hFFB1;
        rom[3][992] = 16'hFFF2;
        rom[3][993] = 16'h0033;
        rom[3][994] = 16'h004F;
        rom[3][995] = 16'h0033;
        rom[3][996] = 16'hFFD5;
        rom[3][997] = 16'hFF9B;
        rom[3][998] = 16'hFF2F;
        rom[3][999] = 16'h003A;
        rom[3][1000] = 16'h0033;
        rom[3][1001] = 16'hFFA9;
        rom[3][1002] = 16'hFF36;
        rom[3][1003] = 16'hFF36;
        rom[3][1004] = 16'hFF9B;
        rom[3][1005] = 16'h0007;
        rom[3][1006] = 16'hFFD5;
        rom[3][1007] = 16'hFED1;
        rom[3][1008] = 16'hFF19;
        rom[3][1009] = 16'hFF7E;
        rom[3][1010] = 16'hFFCD;
        rom[3][1011] = 16'h0007;
        rom[3][1012] = 16'h0000;
        rom[3][1013] = 16'h0000;
        rom[3][1014] = 16'h0000;
        rom[3][1015] = 16'h0000;
        rom[3][1016] = 16'h0000;
        rom[3][1017] = 16'h0000;
        rom[3][1018] = 16'h0000;
        rom[3][1019] = 16'h0000;
        rom[3][1020] = 16'h0000;
        rom[3][1021] = 16'h0000;
        rom[3][1022] = 16'h0000;
        rom[3][1023] = 16'h0000;
        rom[3][1024] = 16'h0000;
        rom[3][1025] = 16'h0000;
        rom[3][1026] = 16'h0000;
        rom[3][1027] = 16'h0000;
        rom[3][1028] = 16'h0000;
        rom[3][1029] = 16'h0000;
        rom[3][1030] = 16'h0000;
        rom[3][1031] = 16'h0000;
        rom[3][1032] = 16'h0000;
        rom[3][1033] = 16'h0000;
        rom[3][1034] = 16'h0000;
        rom[3][1035] = 16'h0000;
        rom[3][1036] = 16'h0000;
        rom[3][1037] = 16'h0000;
        rom[3][1038] = 16'h0000;
        rom[3][1039] = 16'h0000;
        rom[3][1040] = 16'h0000;
        rom[3][1041] = 16'h0000;
        rom[3][1042] = 16'h0000;
        rom[3][1043] = 16'h0000;
        rom[3][1044] = 16'h0000;
        rom[3][1045] = 16'h0000;
        rom[3][1046] = 16'h0000;
        rom[3][1047] = 16'h0000;
        rom[3][1048] = 16'h0000;
        rom[3][1049] = 16'h0000;
        rom[3][1050] = 16'h0000;
        rom[3][1051] = 16'h0000;
        rom[3][1052] = 16'h0000;
        rom[3][1053] = 16'h0000;
        rom[3][1054] = 16'h0000;
        rom[3][1055] = 16'h0000;
        rom[3][1056] = 16'h0000;
        rom[3][1057] = 16'h0000;
        rom[3][1058] = 16'h0000;
        rom[3][1059] = 16'h0000;
        rom[3][1060] = 16'h0000;
        rom[3][1061] = 16'h0000;
        rom[3][1062] = 16'h0000;
        rom[3][1063] = 16'h0000;
        rom[3][1064] = 16'h0000;
        rom[3][1065] = 16'h0000;
        rom[3][1066] = 16'h0000;
        rom[3][1067] = 16'h0000;
        rom[3][1068] = 16'h0000;
        rom[3][1069] = 16'h0000;
        rom[3][1070] = 16'h0000;
        rom[3][1071] = 16'h0000;
        rom[3][1072] = 16'h0000;
        rom[3][1073] = 16'h0000;
        rom[3][1074] = 16'h0000;
        rom[3][1075] = 16'h0000;
        rom[3][1076] = 16'h0000;
        rom[3][1077] = 16'h0000;
        rom[3][1078] = 16'h00E0;
        rom[3][1079] = 16'h0112;
        rom[3][1080] = 16'h00AD;
        rom[3][1081] = 16'h00EE;
        rom[3][1082] = 16'h00AD;
        rom[3][1083] = 16'h00D9;
        rom[3][1084] = 16'h00FD;
        rom[3][1085] = 16'h00EE;
        rom[3][1086] = 16'h00D1;
        rom[3][1087] = 16'h00B4;
        rom[3][1088] = 16'h0082;
        rom[3][1089] = 16'h00A6;
        rom[3][1090] = 16'h009F;
        rom[3][1091] = 16'h00D1;
        rom[3][1092] = 16'h00E7;
        rom[3][1093] = 16'h00A6;
        rom[3][1094] = 16'h0073;
        rom[3][1095] = 16'h0073;
        rom[3][1096] = 16'h0024;
        rom[3][1097] = 16'h015A;
        rom[3][1098] = 16'h01C7;
        rom[3][1099] = 16'h01B1;
        rom[3][1100] = 16'h019B;
        rom[3][1101] = 16'h0169;
        rom[3][1102] = 16'h0121;
        rom[3][1103] = 16'h0170;
        rom[3][1104] = 16'h01DC;
        rom[3][1105] = 16'h00C3;
        rom[3][1106] = 16'h002B;
        rom[3][1107] = 16'h0065;
        rom[3][1108] = 16'h0169;
        rom[3][1109] = 16'h0249;
        rom[3][1110] = 16'h0000;
        rom[3][1111] = 16'h0000;
        rom[3][1112] = 16'h0000;
        rom[3][1113] = 16'h0000;
        rom[3][1114] = 16'h0000;
        rom[3][1115] = 16'h0000;
        rom[3][1116] = 16'h0000;
        rom[3][1117] = 16'h0000;
        rom[3][1118] = 16'h0000;
        rom[3][1119] = 16'h0000;
        rom[3][1120] = 16'h0000;
        rom[3][1121] = 16'h0000;
        rom[3][1122] = 16'h0000;
        rom[3][1123] = 16'h0000;
        rom[3][1124] = 16'h0000;
        rom[3][1125] = 16'h0000;
        rom[3][1126] = 16'h0000;
        rom[3][1127] = 16'h0000;
        rom[3][1128] = 16'h0000;
        rom[3][1129] = 16'h0000;
        rom[3][1130] = 16'h0000;
        rom[3][1131] = 16'h0000;
        rom[3][1132] = 16'h0000;
        rom[3][1133] = 16'h0000;
        rom[3][1134] = 16'h0000;
        rom[3][1135] = 16'h0000;
        rom[3][1136] = 16'h0000;
        rom[3][1137] = 16'h0000;
        rom[3][1138] = 16'h0000;
        rom[3][1139] = 16'h0000;
        rom[3][1140] = 16'h0000;
        rom[3][1141] = 16'h0000;
        rom[3][1142] = 16'h0000;
        rom[3][1143] = 16'h0000;
        rom[3][1144] = 16'h0000;
        rom[3][1145] = 16'h0000;
        rom[3][1146] = 16'h0000;
        rom[3][1147] = 16'h0000;
        rom[3][1148] = 16'h0000;
        rom[3][1149] = 16'h0000;
        rom[3][1150] = 16'h0000;
        rom[3][1151] = 16'h0000;
        rom[3][1152] = 16'h0000;
        rom[3][1153] = 16'h0000;
        rom[3][1154] = 16'h0000;
        rom[3][1155] = 16'h0000;
        rom[3][1156] = 16'h0000;
        rom[3][1157] = 16'h0000;
        rom[3][1158] = 16'h0000;
        rom[3][1159] = 16'h0000;
        rom[3][1160] = 16'h0000;
        rom[3][1161] = 16'h0000;
        rom[3][1162] = 16'h0000;
        rom[3][1163] = 16'h0000;
        rom[3][1164] = 16'h0000;
        rom[3][1165] = 16'h0000;
        rom[3][1166] = 16'h0000;
        rom[3][1167] = 16'h0000;
        rom[3][1168] = 16'h0000;
        rom[3][1169] = 16'h0000;
        rom[3][1170] = 16'h0000;
        rom[3][1171] = 16'h0000;
        rom[3][1172] = 16'h0000;
        rom[3][1173] = 16'h0000;
        rom[3][1174] = 16'h0000;
        rom[3][1175] = 16'h0000;
        rom[3][1176] = 16'hFF5A;
        rom[3][1177] = 16'h0016;
        rom[3][1178] = 16'h0065;
        rom[3][1179] = 16'h005E;
        rom[3][1180] = 16'hFFE3;
        rom[3][1181] = 16'hFF61;
        rom[3][1182] = 16'hFFF9;
        rom[3][1183] = 16'h0048;
        rom[3][1184] = 16'h0041;
        rom[3][1185] = 16'h004F;
        rom[3][1186] = 16'h0024;
        rom[3][1187] = 16'h0041;
        rom[3][1188] = 16'h006C;
        rom[3][1189] = 16'h001D;
        rom[3][1190] = 16'h000E;
        rom[3][1191] = 16'h0065;
        rom[3][1192] = 16'h0065;
        rom[3][1193] = 16'hFFF9;
        rom[3][1194] = 16'hFFBF;
        rom[3][1195] = 16'h003A;
        rom[3][1196] = 16'h005E;
        rom[3][1197] = 16'hFFCD;
        rom[3][1198] = 16'hFFEA;
        rom[3][1199] = 16'h0057;
        rom[3][1200] = 16'h0090;
        rom[3][1201] = 16'h007B;
        rom[3][1202] = 16'h0007;
        rom[3][1203] = 16'hFFDC;
        rom[3][1204] = 16'hFECA;
        rom[3][1205] = 16'hFF27;
        rom[3][1206] = 16'hFFC6;
        rom[3][1207] = 16'hFFB1;
        rom[3][1208] = 16'h0000;
        rom[3][1209] = 16'h0000;
        rom[3][1210] = 16'h0000;
        rom[3][1211] = 16'h0000;
        rom[3][1212] = 16'h0000;
        rom[3][1213] = 16'h0000;
        rom[3][1214] = 16'h0000;
        rom[3][1215] = 16'h0000;
        rom[3][1216] = 16'h0000;
        rom[3][1217] = 16'h0000;
        rom[3][1218] = 16'h0000;
        rom[3][1219] = 16'h0000;
        rom[3][1220] = 16'h0000;
        rom[3][1221] = 16'h0000;
        rom[3][1222] = 16'h0000;
        rom[3][1223] = 16'h0000;
        rom[3][1224] = 16'h0000;
        rom[3][1225] = 16'h0000;
        rom[3][1226] = 16'h0000;
        rom[3][1227] = 16'h0000;
        rom[3][1228] = 16'h0000;
        rom[3][1229] = 16'h0000;
        rom[3][1230] = 16'h0000;
        rom[3][1231] = 16'h0000;
        rom[3][1232] = 16'h0000;
        rom[3][1233] = 16'h0000;
        rom[3][1234] = 16'h0000;
        rom[3][1235] = 16'h0000;
        rom[3][1236] = 16'h0000;
        rom[3][1237] = 16'h0000;
        rom[3][1238] = 16'h0000;
        rom[3][1239] = 16'h0000;
        rom[3][1240] = 16'h0000;
        rom[3][1241] = 16'h0000;
        rom[3][1242] = 16'h0000;
        rom[3][1243] = 16'h0000;
        rom[3][1244] = 16'h0000;
        rom[3][1245] = 16'h0000;
        rom[3][1246] = 16'h0000;
        rom[3][1247] = 16'h0000;
        rom[3][1248] = 16'h0000;
        rom[3][1249] = 16'h0000;
        rom[3][1250] = 16'h0000;
        rom[3][1251] = 16'h0000;
        rom[3][1252] = 16'h0000;
        rom[3][1253] = 16'h0000;
        rom[3][1254] = 16'h0000;
        rom[3][1255] = 16'h0000;
        rom[3][1256] = 16'h0000;
        rom[3][1257] = 16'h0000;
        rom[3][1258] = 16'h0000;
        rom[3][1259] = 16'h0000;
        rom[3][1260] = 16'h0000;
        rom[3][1261] = 16'h0000;
        rom[3][1262] = 16'h0000;
        rom[3][1263] = 16'h0000;
        rom[3][1264] = 16'h0000;
        rom[3][1265] = 16'h0000;
        rom[3][1266] = 16'h0000;
        rom[3][1267] = 16'h0000;
        rom[3][1268] = 16'h0000;
        rom[3][1269] = 16'h0000;
        rom[3][1270] = 16'h0000;
        rom[3][1271] = 16'h0000;
        rom[3][1272] = 16'h0000;
        rom[3][1273] = 16'h0000;
        rom[4][0] = 16'hFF2F;
        rom[4][1] = 16'hFF4C;
        rom[4][2] = 16'hFF4C;
        rom[4][3] = 16'hFF2F;
        rom[4][4] = 16'hFF20;
        rom[4][5] = 16'hFF0B;
        rom[4][6] = 16'hFEF5;
        rom[4][7] = 16'hFEE7;
        rom[4][8] = 16'hFEFC;
        rom[4][9] = 16'hFFA9;
        rom[4][10] = 16'h0000;
        rom[4][11] = 16'h003A;
        rom[4][12] = 16'h004F;
        rom[4][13] = 16'h0024;
        rom[4][14] = 16'hFFB8;
        rom[4][15] = 16'hFF36;
        rom[4][16] = 16'hFEDF;
        rom[4][17] = 16'hFEB4;
        rom[4][18] = 16'hFE9E;
        rom[4][19] = 16'hFE89;
        rom[4][20] = 16'hFE90;
        rom[4][21] = 16'hFE90;
        rom[4][22] = 16'hFE90;
        rom[4][23] = 16'hFE97;
        rom[4][24] = 16'hFEAD;
        rom[4][25] = 16'hFEBB;
        rom[4][26] = 16'hFED8;
        rom[4][27] = 16'hFEE7;
        rom[4][28] = 16'hFEFC;
        rom[4][29] = 16'hFF27;
        rom[4][30] = 16'hFF4C;
        rom[4][31] = 16'hFF5A;
        rom[4][32] = 16'h0000;
        rom[4][33] = 16'h0000;
        rom[4][34] = 16'h0000;
        rom[4][35] = 16'h0000;
        rom[4][36] = 16'h0000;
        rom[4][37] = 16'h0000;
        rom[4][38] = 16'h0000;
        rom[4][39] = 16'h0000;
        rom[4][40] = 16'h0000;
        rom[4][41] = 16'h0000;
        rom[4][42] = 16'h0000;
        rom[4][43] = 16'h0000;
        rom[4][44] = 16'h0000;
        rom[4][45] = 16'h0000;
        rom[4][46] = 16'h0000;
        rom[4][47] = 16'h0000;
        rom[4][48] = 16'h0000;
        rom[4][49] = 16'h0000;
        rom[4][50] = 16'h0000;
        rom[4][51] = 16'h0000;
        rom[4][52] = 16'h0000;
        rom[4][53] = 16'h0000;
        rom[4][54] = 16'h0000;
        rom[4][55] = 16'h0000;
        rom[4][56] = 16'h0000;
        rom[4][57] = 16'h0000;
        rom[4][58] = 16'h0000;
        rom[4][59] = 16'h0000;
        rom[4][60] = 16'h0000;
        rom[4][61] = 16'h0000;
        rom[4][62] = 16'h0000;
        rom[4][63] = 16'h0000;
        rom[4][64] = 16'h0000;
        rom[4][65] = 16'h0000;
        rom[4][66] = 16'h0000;
        rom[4][67] = 16'h0000;
        rom[4][68] = 16'h0000;
        rom[4][69] = 16'h0000;
        rom[4][70] = 16'h0000;
        rom[4][71] = 16'h0000;
        rom[4][72] = 16'h0000;
        rom[4][73] = 16'h0000;
        rom[4][74] = 16'h0000;
        rom[4][75] = 16'h0000;
        rom[4][76] = 16'h0000;
        rom[4][77] = 16'h0000;
        rom[4][78] = 16'h0000;
        rom[4][79] = 16'h0000;
        rom[4][80] = 16'h0000;
        rom[4][81] = 16'h0000;
        rom[4][82] = 16'h0000;
        rom[4][83] = 16'h0000;
        rom[4][84] = 16'h0000;
        rom[4][85] = 16'h0000;
        rom[4][86] = 16'h0000;
        rom[4][87] = 16'h0000;
        rom[4][88] = 16'h0000;
        rom[4][89] = 16'h0000;
        rom[4][90] = 16'h0000;
        rom[4][91] = 16'h0000;
        rom[4][92] = 16'h0000;
        rom[4][93] = 16'h0000;
        rom[4][94] = 16'h0000;
        rom[4][95] = 16'h0000;
        rom[4][96] = 16'h0000;
        rom[4][97] = 16'h0000;
        rom[4][98] = 16'h0098;
        rom[4][99] = 16'h0082;
        rom[4][100] = 16'h005E;
        rom[4][101] = 16'h0048;
        rom[4][102] = 16'h0024;
        rom[4][103] = 16'hFFE3;
        rom[4][104] = 16'hFFBF;
        rom[4][105] = 16'hFFC6;
        rom[4][106] = 16'h0000;
        rom[4][107] = 16'h0048;
        rom[4][108] = 16'h001D;
        rom[4][109] = 16'h001D;
        rom[4][110] = 16'h0024;
        rom[4][111] = 16'h0033;
        rom[4][112] = 16'h0041;
        rom[4][113] = 16'h004F;
        rom[4][114] = 16'h0016;
        rom[4][115] = 16'hFFE3;
        rom[4][116] = 16'hFFEA;
        rom[4][117] = 16'hFFB1;
        rom[4][118] = 16'hFF7E;
        rom[4][119] = 16'hFF94;
        rom[4][120] = 16'hFFA9;
        rom[4][121] = 16'hFFA2;
        rom[4][122] = 16'hFFB1;
        rom[4][123] = 16'hFFC6;
        rom[4][124] = 16'hFFD5;
        rom[4][125] = 16'hFFE3;
        rom[4][126] = 16'hFFEA;
        rom[4][127] = 16'h0024;
        rom[4][128] = 16'h0057;
        rom[4][129] = 16'h009F;
        rom[4][130] = 16'h0000;
        rom[4][131] = 16'h0000;
        rom[4][132] = 16'h0000;
        rom[4][133] = 16'h0000;
        rom[4][134] = 16'h0000;
        rom[4][135] = 16'h0000;
        rom[4][136] = 16'h0000;
        rom[4][137] = 16'h0000;
        rom[4][138] = 16'h0000;
        rom[4][139] = 16'h0000;
        rom[4][140] = 16'h0000;
        rom[4][141] = 16'h0000;
        rom[4][142] = 16'h0000;
        rom[4][143] = 16'h0000;
        rom[4][144] = 16'h0000;
        rom[4][145] = 16'h0000;
        rom[4][146] = 16'h0000;
        rom[4][147] = 16'h0000;
        rom[4][148] = 16'h0000;
        rom[4][149] = 16'h0000;
        rom[4][150] = 16'h0000;
        rom[4][151] = 16'h0000;
        rom[4][152] = 16'h0000;
        rom[4][153] = 16'h0000;
        rom[4][154] = 16'h0000;
        rom[4][155] = 16'h0000;
        rom[4][156] = 16'h0000;
        rom[4][157] = 16'h0000;
        rom[4][158] = 16'h0000;
        rom[4][159] = 16'h0000;
        rom[4][160] = 16'h0000;
        rom[4][161] = 16'h0000;
        rom[4][162] = 16'h0000;
        rom[4][163] = 16'h0000;
        rom[4][164] = 16'h0000;
        rom[4][165] = 16'h0000;
        rom[4][166] = 16'h0000;
        rom[4][167] = 16'h0000;
        rom[4][168] = 16'h0000;
        rom[4][169] = 16'h0000;
        rom[4][170] = 16'h0000;
        rom[4][171] = 16'h0000;
        rom[4][172] = 16'h0000;
        rom[4][173] = 16'h0000;
        rom[4][174] = 16'h0000;
        rom[4][175] = 16'h0000;
        rom[4][176] = 16'h0000;
        rom[4][177] = 16'h0000;
        rom[4][178] = 16'h0000;
        rom[4][179] = 16'h0000;
        rom[4][180] = 16'h0000;
        rom[4][181] = 16'h0000;
        rom[4][182] = 16'h0000;
        rom[4][183] = 16'h0000;
        rom[4][184] = 16'h0000;
        rom[4][185] = 16'h0000;
        rom[4][186] = 16'h0000;
        rom[4][187] = 16'h0000;
        rom[4][188] = 16'h0000;
        rom[4][189] = 16'h0000;
        rom[4][190] = 16'h0000;
        rom[4][191] = 16'h0000;
        rom[4][192] = 16'h0000;
        rom[4][193] = 16'h0000;
        rom[4][194] = 16'h0000;
        rom[4][195] = 16'h0000;
        rom[4][196] = 16'hFF77;
        rom[4][197] = 16'hFF2F;
        rom[4][198] = 16'hFF27;
        rom[4][199] = 16'hFF7E;
        rom[4][200] = 16'hFF94;
        rom[4][201] = 16'hFF70;
        rom[4][202] = 16'hFF68;
        rom[4][203] = 16'hFF94;
        rom[4][204] = 16'hFFB1;
        rom[4][205] = 16'hFF85;
        rom[4][206] = 16'hFF9B;
        rom[4][207] = 16'hFF70;
        rom[4][208] = 16'hFF19;
        rom[4][209] = 16'hFF20;
        rom[4][210] = 16'hFF4C;
        rom[4][211] = 16'hFF7E;
        rom[4][212] = 16'hFFA2;
        rom[4][213] = 16'hFFF2;
        rom[4][214] = 16'h0057;
        rom[4][215] = 16'h005E;
        rom[4][216] = 16'h0048;
        rom[4][217] = 16'h0033;
        rom[4][218] = 16'h001D;
        rom[4][219] = 16'hFFF9;
        rom[4][220] = 16'hFFB1;
        rom[4][221] = 16'hFF9B;
        rom[4][222] = 16'hFFB1;
        rom[4][223] = 16'hFFBF;
        rom[4][224] = 16'hFFB8;
        rom[4][225] = 16'hFFA2;
        rom[4][226] = 16'hFFC6;
        rom[4][227] = 16'hFFEA;
        rom[4][228] = 16'h0000;
        rom[4][229] = 16'h0000;
        rom[4][230] = 16'h0000;
        rom[4][231] = 16'h0000;
        rom[4][232] = 16'h0000;
        rom[4][233] = 16'h0000;
        rom[4][234] = 16'h0000;
        rom[4][235] = 16'h0000;
        rom[4][236] = 16'h0000;
        rom[4][237] = 16'h0000;
        rom[4][238] = 16'h0000;
        rom[4][239] = 16'h0000;
        rom[4][240] = 16'h0000;
        rom[4][241] = 16'h0000;
        rom[4][242] = 16'h0000;
        rom[4][243] = 16'h0000;
        rom[4][244] = 16'h0000;
        rom[4][245] = 16'h0000;
        rom[4][246] = 16'h0000;
        rom[4][247] = 16'h0000;
        rom[4][248] = 16'h0000;
        rom[4][249] = 16'h0000;
        rom[4][250] = 16'h0000;
        rom[4][251] = 16'h0000;
        rom[4][252] = 16'h0000;
        rom[4][253] = 16'h0000;
        rom[4][254] = 16'h0000;
        rom[4][255] = 16'h0000;
        rom[4][256] = 16'h0000;
        rom[4][257] = 16'h0000;
        rom[4][258] = 16'h0000;
        rom[4][259] = 16'h0000;
        rom[4][260] = 16'h0000;
        rom[4][261] = 16'h0000;
        rom[4][262] = 16'h0000;
        rom[4][263] = 16'h0000;
        rom[4][264] = 16'h0000;
        rom[4][265] = 16'h0000;
        rom[4][266] = 16'h0000;
        rom[4][267] = 16'h0000;
        rom[4][268] = 16'h0000;
        rom[4][269] = 16'h0000;
        rom[4][270] = 16'h0000;
        rom[4][271] = 16'h0000;
        rom[4][272] = 16'h0000;
        rom[4][273] = 16'h0000;
        rom[4][274] = 16'h0000;
        rom[4][275] = 16'h0000;
        rom[4][276] = 16'h0000;
        rom[4][277] = 16'h0000;
        rom[4][278] = 16'h0000;
        rom[4][279] = 16'h0000;
        rom[4][280] = 16'h0000;
        rom[4][281] = 16'h0000;
        rom[4][282] = 16'h0000;
        rom[4][283] = 16'h0000;
        rom[4][284] = 16'h0000;
        rom[4][285] = 16'h0000;
        rom[4][286] = 16'h0000;
        rom[4][287] = 16'h0000;
        rom[4][288] = 16'h0000;
        rom[4][289] = 16'h0000;
        rom[4][290] = 16'h0000;
        rom[4][291] = 16'h0000;
        rom[4][292] = 16'h0000;
        rom[4][293] = 16'h0000;
        rom[4][294] = 16'hFFF2;
        rom[4][295] = 16'hFF77;
        rom[4][296] = 16'hFF3D;
        rom[4][297] = 16'hFFA9;
        rom[4][298] = 16'hFFEA;
        rom[4][299] = 16'hFFF2;
        rom[4][300] = 16'hFF70;
        rom[4][301] = 16'hFF19;
        rom[4][302] = 16'hFEEE;
        rom[4][303] = 16'hFED8;
        rom[4][304] = 16'hFE73;
        rom[4][305] = 16'hFE0E;
        rom[4][306] = 16'hFE2B;
        rom[4][307] = 16'hFE90;
        rom[4][308] = 16'hFED8;
        rom[4][309] = 16'hFEBB;
        rom[4][310] = 16'hFF27;
        rom[4][311] = 16'hFFCD;
        rom[4][312] = 16'h007B;
        rom[4][313] = 16'h007B;
        rom[4][314] = 16'h0048;
        rom[4][315] = 16'h0033;
        rom[4][316] = 16'h002B;
        rom[4][317] = 16'h003A;
        rom[4][318] = 16'h0007;
        rom[4][319] = 16'hFFC6;
        rom[4][320] = 16'hFFD5;
        rom[4][321] = 16'hFFC6;
        rom[4][322] = 16'hFF77;
        rom[4][323] = 16'hFFB8;
        rom[4][324] = 16'h001D;
        rom[4][325] = 16'h0033;
        rom[4][326] = 16'h0000;
        rom[4][327] = 16'h0000;
        rom[4][328] = 16'h0000;
        rom[4][329] = 16'h0000;
        rom[4][330] = 16'h0000;
        rom[4][331] = 16'h0000;
        rom[4][332] = 16'h0000;
        rom[4][333] = 16'h0000;
        rom[4][334] = 16'h0000;
        rom[4][335] = 16'h0000;
        rom[4][336] = 16'h0000;
        rom[4][337] = 16'h0000;
        rom[4][338] = 16'h0000;
        rom[4][339] = 16'h0000;
        rom[4][340] = 16'h0000;
        rom[4][341] = 16'h0000;
        rom[4][342] = 16'h0000;
        rom[4][343] = 16'h0000;
        rom[4][344] = 16'h0000;
        rom[4][345] = 16'h0000;
        rom[4][346] = 16'h0000;
        rom[4][347] = 16'h0000;
        rom[4][348] = 16'h0000;
        rom[4][349] = 16'h0000;
        rom[4][350] = 16'h0000;
        rom[4][351] = 16'h0000;
        rom[4][352] = 16'h0000;
        rom[4][353] = 16'h0000;
        rom[4][354] = 16'h0000;
        rom[4][355] = 16'h0000;
        rom[4][356] = 16'h0000;
        rom[4][357] = 16'h0000;
        rom[4][358] = 16'h0000;
        rom[4][359] = 16'h0000;
        rom[4][360] = 16'h0000;
        rom[4][361] = 16'h0000;
        rom[4][362] = 16'h0000;
        rom[4][363] = 16'h0000;
        rom[4][364] = 16'h0000;
        rom[4][365] = 16'h0000;
        rom[4][366] = 16'h0000;
        rom[4][367] = 16'h0000;
        rom[4][368] = 16'h0000;
        rom[4][369] = 16'h0000;
        rom[4][370] = 16'h0000;
        rom[4][371] = 16'h0000;
        rom[4][372] = 16'h0000;
        rom[4][373] = 16'h0000;
        rom[4][374] = 16'h0000;
        rom[4][375] = 16'h0000;
        rom[4][376] = 16'h0000;
        rom[4][377] = 16'h0000;
        rom[4][378] = 16'h0000;
        rom[4][379] = 16'h0000;
        rom[4][380] = 16'h0000;
        rom[4][381] = 16'h0000;
        rom[4][382] = 16'h0000;
        rom[4][383] = 16'h0000;
        rom[4][384] = 16'h0000;
        rom[4][385] = 16'h0000;
        rom[4][386] = 16'h0000;
        rom[4][387] = 16'h0000;
        rom[4][388] = 16'h0000;
        rom[4][389] = 16'h0000;
        rom[4][390] = 16'h0000;
        rom[4][391] = 16'h0000;
        rom[4][392] = 16'h0057;
        rom[4][393] = 16'hFFDC;
        rom[4][394] = 16'hFF77;
        rom[4][395] = 16'hFF70;
        rom[4][396] = 16'hFFCD;
        rom[4][397] = 16'h0024;
        rom[4][398] = 16'hFFF2;
        rom[4][399] = 16'hFFA2;
        rom[4][400] = 16'hFFF9;
        rom[4][401] = 16'hFEBB;
        rom[4][402] = 16'hFE81;
        rom[4][403] = 16'hFE39;
        rom[4][404] = 16'hFE00;
        rom[4][405] = 16'hFE0E;
        rom[4][406] = 16'hFE41;
        rom[4][407] = 16'hFF36;
        rom[4][408] = 16'h002B;
        rom[4][409] = 16'h005E;
        rom[4][410] = 16'h0073;
        rom[4][411] = 16'h00C3;
        rom[4][412] = 16'h00A6;
        rom[4][413] = 16'h0082;
        rom[4][414] = 16'h007B;
        rom[4][415] = 16'h004F;
        rom[4][416] = 16'h0033;
        rom[4][417] = 16'h0041;
        rom[4][418] = 16'h0041;
        rom[4][419] = 16'hFFF2;
        rom[4][420] = 16'hFF77;
        rom[4][421] = 16'hFF94;
        rom[4][422] = 16'h002B;
        rom[4][423] = 16'h00D9;
        rom[4][424] = 16'h0000;
        rom[4][425] = 16'h0000;
        rom[4][426] = 16'h0000;
        rom[4][427] = 16'h0000;
        rom[4][428] = 16'h0000;
        rom[4][429] = 16'h0000;
        rom[4][430] = 16'h0000;
        rom[4][431] = 16'h0000;
        rom[4][432] = 16'h0000;
        rom[4][433] = 16'h0000;
        rom[4][434] = 16'h0000;
        rom[4][435] = 16'h0000;
        rom[4][436] = 16'h0000;
        rom[4][437] = 16'h0000;
        rom[4][438] = 16'h0000;
        rom[4][439] = 16'h0000;
        rom[4][440] = 16'h0000;
        rom[4][441] = 16'h0000;
        rom[4][442] = 16'h0000;
        rom[4][443] = 16'h0000;
        rom[4][444] = 16'h0000;
        rom[4][445] = 16'h0000;
        rom[4][446] = 16'h0000;
        rom[4][447] = 16'h0000;
        rom[4][448] = 16'h0000;
        rom[4][449] = 16'h0000;
        rom[4][450] = 16'h0000;
        rom[4][451] = 16'h0000;
        rom[4][452] = 16'h0000;
        rom[4][453] = 16'h0000;
        rom[4][454] = 16'h0000;
        rom[4][455] = 16'h0000;
        rom[4][456] = 16'h0000;
        rom[4][457] = 16'h0000;
        rom[4][458] = 16'h0000;
        rom[4][459] = 16'h0000;
        rom[4][460] = 16'h0000;
        rom[4][461] = 16'h0000;
        rom[4][462] = 16'h0000;
        rom[4][463] = 16'h0000;
        rom[4][464] = 16'h0000;
        rom[4][465] = 16'h0000;
        rom[4][466] = 16'h0000;
        rom[4][467] = 16'h0000;
        rom[4][468] = 16'h0000;
        rom[4][469] = 16'h0000;
        rom[4][470] = 16'h0000;
        rom[4][471] = 16'h0000;
        rom[4][472] = 16'h0000;
        rom[4][473] = 16'h0000;
        rom[4][474] = 16'h0000;
        rom[4][475] = 16'h0000;
        rom[4][476] = 16'h0000;
        rom[4][477] = 16'h0000;
        rom[4][478] = 16'h0000;
        rom[4][479] = 16'h0000;
        rom[4][480] = 16'h0000;
        rom[4][481] = 16'h0000;
        rom[4][482] = 16'h0000;
        rom[4][483] = 16'h0000;
        rom[4][484] = 16'h0000;
        rom[4][485] = 16'h0000;
        rom[4][486] = 16'h0000;
        rom[4][487] = 16'h0000;
        rom[4][488] = 16'h0000;
        rom[4][489] = 16'h0000;
        rom[4][490] = 16'hFFD5;
        rom[4][491] = 16'h006C;
        rom[4][492] = 16'h0065;
        rom[4][493] = 16'hFFEA;
        rom[4][494] = 16'hFF9B;
        rom[4][495] = 16'hFFCD;
        rom[4][496] = 16'h0024;
        rom[4][497] = 16'h006C;
        rom[4][498] = 16'h00AD;
        rom[4][499] = 16'h01F2;
        rom[4][500] = 16'h0225;
        rom[4][501] = 16'h019B;
        rom[4][502] = 16'h013E;
        rom[4][503] = 16'h0136;
        rom[4][504] = 16'h00D9;
        rom[4][505] = 16'h009F;
        rom[4][506] = 16'h00EE;
        rom[4][507] = 16'h00BC;
        rom[4][508] = 16'h0048;
        rom[4][509] = 16'h0090;
        rom[4][510] = 16'h0089;
        rom[4][511] = 16'h0082;
        rom[4][512] = 16'h001D;
        rom[4][513] = 16'hFFBF;
        rom[4][514] = 16'hFFC6;
        rom[4][515] = 16'h0016;
        rom[4][516] = 16'h004F;
        rom[4][517] = 16'hFFF9;
        rom[4][518] = 16'hFFBF;
        rom[4][519] = 16'hFF9B;
        rom[4][520] = 16'h0000;
        rom[4][521] = 16'h003A;
        rom[4][522] = 16'h0000;
        rom[4][523] = 16'h0000;
        rom[4][524] = 16'h0000;
        rom[4][525] = 16'h0000;
        rom[4][526] = 16'h0000;
        rom[4][527] = 16'h0000;
        rom[4][528] = 16'h0000;
        rom[4][529] = 16'h0000;
        rom[4][530] = 16'h0000;
        rom[4][531] = 16'h0000;
        rom[4][532] = 16'h0000;
        rom[4][533] = 16'h0000;
        rom[4][534] = 16'h0000;
        rom[4][535] = 16'h0000;
        rom[4][536] = 16'h0000;
        rom[4][537] = 16'h0000;
        rom[4][538] = 16'h0000;
        rom[4][539] = 16'h0000;
        rom[4][540] = 16'h0000;
        rom[4][541] = 16'h0000;
        rom[4][542] = 16'h0000;
        rom[4][543] = 16'h0000;
        rom[4][544] = 16'h0000;
        rom[4][545] = 16'h0000;
        rom[4][546] = 16'h0000;
        rom[4][547] = 16'h0000;
        rom[4][548] = 16'h0000;
        rom[4][549] = 16'h0000;
        rom[4][550] = 16'h0000;
        rom[4][551] = 16'h0000;
        rom[4][552] = 16'h0000;
        rom[4][553] = 16'h0000;
        rom[4][554] = 16'h0000;
        rom[4][555] = 16'h0000;
        rom[4][556] = 16'h0000;
        rom[4][557] = 16'h0000;
        rom[4][558] = 16'h0000;
        rom[4][559] = 16'h0000;
        rom[4][560] = 16'h0000;
        rom[4][561] = 16'h0000;
        rom[4][562] = 16'h0000;
        rom[4][563] = 16'h0000;
        rom[4][564] = 16'h0000;
        rom[4][565] = 16'h0000;
        rom[4][566] = 16'h0000;
        rom[4][567] = 16'h0000;
        rom[4][568] = 16'h0000;
        rom[4][569] = 16'h0000;
        rom[4][570] = 16'h0000;
        rom[4][571] = 16'h0000;
        rom[4][572] = 16'h0000;
        rom[4][573] = 16'h0000;
        rom[4][574] = 16'h0000;
        rom[4][575] = 16'h0000;
        rom[4][576] = 16'h0000;
        rom[4][577] = 16'h0000;
        rom[4][578] = 16'h0000;
        rom[4][579] = 16'h0000;
        rom[4][580] = 16'h0000;
        rom[4][581] = 16'h0000;
        rom[4][582] = 16'h0000;
        rom[4][583] = 16'h0000;
        rom[4][584] = 16'h0000;
        rom[4][585] = 16'h0000;
        rom[4][586] = 16'h0000;
        rom[4][587] = 16'h0000;
        rom[4][588] = 16'h0007;
        rom[4][589] = 16'h0033;
        rom[4][590] = 16'h0024;
        rom[4][591] = 16'h001D;
        rom[4][592] = 16'h0065;
        rom[4][593] = 16'h0073;
        rom[4][594] = 16'h004F;
        rom[4][595] = 16'h00A6;
        rom[4][596] = 16'h007B;
        rom[4][597] = 16'hFFD5;
        rom[4][598] = 16'hFFBF;
        rom[4][599] = 16'hFF94;
        rom[4][600] = 16'hFFA9;
        rom[4][601] = 16'hFFEA;
        rom[4][602] = 16'h0000;
        rom[4][603] = 16'hFFA2;
        rom[4][604] = 16'hFFF9;
        rom[4][605] = 16'h000E;
        rom[4][606] = 16'h0024;
        rom[4][607] = 16'h0057;
        rom[4][608] = 16'hFFA2;
        rom[4][609] = 16'hFF9B;
        rom[4][610] = 16'hFFE3;
        rom[4][611] = 16'hFFDC;
        rom[4][612] = 16'hFFDC;
        rom[4][613] = 16'h0007;
        rom[4][614] = 16'h005E;
        rom[4][615] = 16'h0033;
        rom[4][616] = 16'h0065;
        rom[4][617] = 16'h0082;
        rom[4][618] = 16'hFFD5;
        rom[4][619] = 16'hFF27;
        rom[4][620] = 16'h0000;
        rom[4][621] = 16'h0000;
        rom[4][622] = 16'h0000;
        rom[4][623] = 16'h0000;
        rom[4][624] = 16'h0000;
        rom[4][625] = 16'h0000;
        rom[4][626] = 16'h0000;
        rom[4][627] = 16'h0000;
        rom[4][628] = 16'h0000;
        rom[4][629] = 16'h0000;
        rom[4][630] = 16'h0000;
        rom[4][631] = 16'h0000;
        rom[4][632] = 16'h0000;
        rom[4][633] = 16'h0000;
        rom[4][634] = 16'h0000;
        rom[4][635] = 16'h0000;
        rom[4][636] = 16'h0000;
        rom[4][637] = 16'h0000;
        rom[4][638] = 16'h0000;
        rom[4][639] = 16'h0000;
        rom[4][640] = 16'h0000;
        rom[4][641] = 16'h0000;
        rom[4][642] = 16'h0000;
        rom[4][643] = 16'h0000;
        rom[4][644] = 16'h0000;
        rom[4][645] = 16'h0000;
        rom[4][646] = 16'h0000;
        rom[4][647] = 16'h0000;
        rom[4][648] = 16'h0000;
        rom[4][649] = 16'h0000;
        rom[4][650] = 16'h0000;
        rom[4][651] = 16'h0000;
        rom[4][652] = 16'h0000;
        rom[4][653] = 16'h0000;
        rom[4][654] = 16'h0000;
        rom[4][655] = 16'h0000;
        rom[4][656] = 16'h0000;
        rom[4][657] = 16'h0000;
        rom[4][658] = 16'h0000;
        rom[4][659] = 16'h0000;
        rom[4][660] = 16'h0000;
        rom[4][661] = 16'h0000;
        rom[4][662] = 16'h0000;
        rom[4][663] = 16'h0000;
        rom[4][664] = 16'h0000;
        rom[4][665] = 16'h0000;
        rom[4][666] = 16'h0000;
        rom[4][667] = 16'h0000;
        rom[4][668] = 16'h0000;
        rom[4][669] = 16'h0000;
        rom[4][670] = 16'h0000;
        rom[4][671] = 16'h0000;
        rom[4][672] = 16'h0000;
        rom[4][673] = 16'h0000;
        rom[4][674] = 16'h0000;
        rom[4][675] = 16'h0000;
        rom[4][676] = 16'h0000;
        rom[4][677] = 16'h0000;
        rom[4][678] = 16'h0000;
        rom[4][679] = 16'h0000;
        rom[4][680] = 16'h0000;
        rom[4][681] = 16'h0000;
        rom[4][682] = 16'h0000;
        rom[4][683] = 16'h0000;
        rom[4][684] = 16'h0000;
        rom[4][685] = 16'h0000;
        rom[4][686] = 16'hFFA2;
        rom[4][687] = 16'hFF27;
        rom[4][688] = 16'hFEFC;
        rom[4][689] = 16'hFF77;
        rom[4][690] = 16'hFF9B;
        rom[4][691] = 16'hFFA9;
        rom[4][692] = 16'hFFDC;
        rom[4][693] = 16'h004F;
        rom[4][694] = 16'hFFC6;
        rom[4][695] = 16'hFED1;
        rom[4][696] = 16'hFED8;
        rom[4][697] = 16'hFECA;
        rom[4][698] = 16'hFED8;
        rom[4][699] = 16'hFF03;
        rom[4][700] = 16'hFEFC;
        rom[4][701] = 16'hFF44;
        rom[4][702] = 16'hFFF2;
        rom[4][703] = 16'h000E;
        rom[4][704] = 16'h005E;
        rom[4][705] = 16'h00B4;
        rom[4][706] = 16'hFFA9;
        rom[4][707] = 16'hFF0B;
        rom[4][708] = 16'hFFB8;
        rom[4][709] = 16'h0000;
        rom[4][710] = 16'hFF94;
        rom[4][711] = 16'hFF7E;
        rom[4][712] = 16'hFFA9;
        rom[4][713] = 16'hFFC6;
        rom[4][714] = 16'hFFB1;
        rom[4][715] = 16'hFFC6;
        rom[4][716] = 16'hFFA9;
        rom[4][717] = 16'hFF12;
        rom[4][718] = 16'h0000;
        rom[4][719] = 16'h0000;
        rom[4][720] = 16'h0000;
        rom[4][721] = 16'h0000;
        rom[4][722] = 16'h0000;
        rom[4][723] = 16'h0000;
        rom[4][724] = 16'h0000;
        rom[4][725] = 16'h0000;
        rom[4][726] = 16'h0000;
        rom[4][727] = 16'h0000;
        rom[4][728] = 16'h0000;
        rom[4][729] = 16'h0000;
        rom[4][730] = 16'h0000;
        rom[4][731] = 16'h0000;
        rom[4][732] = 16'h0000;
        rom[4][733] = 16'h0000;
        rom[4][734] = 16'h0000;
        rom[4][735] = 16'h0000;
        rom[4][736] = 16'h0000;
        rom[4][737] = 16'h0000;
        rom[4][738] = 16'h0000;
        rom[4][739] = 16'h0000;
        rom[4][740] = 16'h0000;
        rom[4][741] = 16'h0000;
        rom[4][742] = 16'h0000;
        rom[4][743] = 16'h0000;
        rom[4][744] = 16'h0000;
        rom[4][745] = 16'h0000;
        rom[4][746] = 16'h0000;
        rom[4][747] = 16'h0000;
        rom[4][748] = 16'h0000;
        rom[4][749] = 16'h0000;
        rom[4][750] = 16'h0000;
        rom[4][751] = 16'h0000;
        rom[4][752] = 16'h0000;
        rom[4][753] = 16'h0000;
        rom[4][754] = 16'h0000;
        rom[4][755] = 16'h0000;
        rom[4][756] = 16'h0000;
        rom[4][757] = 16'h0000;
        rom[4][758] = 16'h0000;
        rom[4][759] = 16'h0000;
        rom[4][760] = 16'h0000;
        rom[4][761] = 16'h0000;
        rom[4][762] = 16'h0000;
        rom[4][763] = 16'h0000;
        rom[4][764] = 16'h0000;
        rom[4][765] = 16'h0000;
        rom[4][766] = 16'h0000;
        rom[4][767] = 16'h0000;
        rom[4][768] = 16'h0000;
        rom[4][769] = 16'h0000;
        rom[4][770] = 16'h0000;
        rom[4][771] = 16'h0000;
        rom[4][772] = 16'h0000;
        rom[4][773] = 16'h0000;
        rom[4][774] = 16'h0000;
        rom[4][775] = 16'h0000;
        rom[4][776] = 16'h0000;
        rom[4][777] = 16'h0000;
        rom[4][778] = 16'h0000;
        rom[4][779] = 16'h0000;
        rom[4][780] = 16'h0000;
        rom[4][781] = 16'h0000;
        rom[4][782] = 16'h0000;
        rom[4][783] = 16'h0000;
        rom[4][784] = 16'hFE39;
        rom[4][785] = 16'hFDDB;
        rom[4][786] = 16'hFE0E;
        rom[4][787] = 16'hFEC2;
        rom[4][788] = 16'hFE0E;
        rom[4][789] = 16'hFD93;
        rom[4][790] = 16'hFE07;
        rom[4][791] = 16'hFECA;
        rom[4][792] = 16'hFE39;
        rom[4][793] = 16'hFD20;
        rom[4][794] = 16'hFCB4;
        rom[4][795] = 16'hFCFC;
        rom[4][796] = 16'hFD19;
        rom[4][797] = 16'hFCE6;
        rom[4][798] = 16'hFCD8;
        rom[4][799] = 16'hFD8C;
        rom[4][800] = 16'hFE56;
        rom[4][801] = 16'hFEDF;
        rom[4][802] = 16'hFF3D;
        rom[4][803] = 16'hFEF5;
        rom[4][804] = 16'hFE32;
        rom[4][805] = 16'hFDB0;
        rom[4][806] = 16'hFE00;
        rom[4][807] = 16'hFE65;
        rom[4][808] = 16'hFE65;
        rom[4][809] = 16'hFE1C;
        rom[4][810] = 16'hFDCD;
        rom[4][811] = 16'hFE7A;
        rom[4][812] = 16'hFE1C;
        rom[4][813] = 16'hFD5A;
        rom[4][814] = 16'hFD19;
        rom[4][815] = 16'hFDC6;
        rom[4][816] = 16'h0000;
        rom[4][817] = 16'h0000;
        rom[4][818] = 16'h0000;
        rom[4][819] = 16'h0000;
        rom[4][820] = 16'h0000;
        rom[4][821] = 16'h0000;
        rom[4][822] = 16'h0000;
        rom[4][823] = 16'h0000;
        rom[4][824] = 16'h0000;
        rom[4][825] = 16'h0000;
        rom[4][826] = 16'h0000;
        rom[4][827] = 16'h0000;
        rom[4][828] = 16'h0000;
        rom[4][829] = 16'h0000;
        rom[4][830] = 16'h0000;
        rom[4][831] = 16'h0000;
        rom[4][832] = 16'h0000;
        rom[4][833] = 16'h0000;
        rom[4][834] = 16'h0000;
        rom[4][835] = 16'h0000;
        rom[4][836] = 16'h0000;
        rom[4][837] = 16'h0000;
        rom[4][838] = 16'h0000;
        rom[4][839] = 16'h0000;
        rom[4][840] = 16'h0000;
        rom[4][841] = 16'h0000;
        rom[4][842] = 16'h0000;
        rom[4][843] = 16'h0000;
        rom[4][844] = 16'h0000;
        rom[4][845] = 16'h0000;
        rom[4][846] = 16'h0000;
        rom[4][847] = 16'h0000;
        rom[4][848] = 16'h0000;
        rom[4][849] = 16'h0000;
        rom[4][850] = 16'h0000;
        rom[4][851] = 16'h0000;
        rom[4][852] = 16'h0000;
        rom[4][853] = 16'h0000;
        rom[4][854] = 16'h0000;
        rom[4][855] = 16'h0000;
        rom[4][856] = 16'h0000;
        rom[4][857] = 16'h0000;
        rom[4][858] = 16'h0000;
        rom[4][859] = 16'h0000;
        rom[4][860] = 16'h0000;
        rom[4][861] = 16'h0000;
        rom[4][862] = 16'h0000;
        rom[4][863] = 16'h0000;
        rom[4][864] = 16'h0000;
        rom[4][865] = 16'h0000;
        rom[4][866] = 16'h0000;
        rom[4][867] = 16'h0000;
        rom[4][868] = 16'h0000;
        rom[4][869] = 16'h0000;
        rom[4][870] = 16'h0000;
        rom[4][871] = 16'h0000;
        rom[4][872] = 16'h0000;
        rom[4][873] = 16'h0000;
        rom[4][874] = 16'h0000;
        rom[4][875] = 16'h0000;
        rom[4][876] = 16'h0000;
        rom[4][877] = 16'h0000;
        rom[4][878] = 16'h0000;
        rom[4][879] = 16'h0000;
        rom[4][880] = 16'h0000;
        rom[4][881] = 16'h0000;
        rom[4][882] = 16'hFEFC;
        rom[4][883] = 16'hFEC2;
        rom[4][884] = 16'hFEAD;
        rom[4][885] = 16'hFEFC;
        rom[4][886] = 16'hFF20;
        rom[4][887] = 16'hFECA;
        rom[4][888] = 16'hFEE7;
        rom[4][889] = 16'hFF4C;
        rom[4][890] = 16'hFF61;
        rom[4][891] = 16'hFFE3;
        rom[4][892] = 16'h00EE;
        rom[4][893] = 16'h01B1;
        rom[4][894] = 16'h0177;
        rom[4][895] = 16'h00C3;
        rom[4][896] = 16'hFFC6;
        rom[4][897] = 16'hFFB8;
        rom[4][898] = 16'h004F;
        rom[4][899] = 16'h0136;
        rom[4][900] = 16'h007B;
        rom[4][901] = 16'hFFDC;
        rom[4][902] = 16'hFFB1;
        rom[4][903] = 16'hFF44;
        rom[4][904] = 16'hFF19;
        rom[4][905] = 16'hFED8;
        rom[4][906] = 16'hFEE7;
        rom[4][907] = 16'hFEEE;
        rom[4][908] = 16'hFF27;
        rom[4][909] = 16'hFF61;
        rom[4][910] = 16'hFF94;
        rom[4][911] = 16'hFEFC;
        rom[4][912] = 16'hFE65;
        rom[4][913] = 16'hFED8;
        rom[4][914] = 16'h0000;
        rom[4][915] = 16'h0000;
        rom[4][916] = 16'h0000;
        rom[4][917] = 16'h0000;
        rom[4][918] = 16'h0000;
        rom[4][919] = 16'h0000;
        rom[4][920] = 16'h0000;
        rom[4][921] = 16'h0000;
        rom[4][922] = 16'h0000;
        rom[4][923] = 16'h0000;
        rom[4][924] = 16'h0000;
        rom[4][925] = 16'h0000;
        rom[4][926] = 16'h0000;
        rom[4][927] = 16'h0000;
        rom[4][928] = 16'h0000;
        rom[4][929] = 16'h0000;
        rom[4][930] = 16'h0000;
        rom[4][931] = 16'h0000;
        rom[4][932] = 16'h0000;
        rom[4][933] = 16'h0000;
        rom[4][934] = 16'h0000;
        rom[4][935] = 16'h0000;
        rom[4][936] = 16'h0000;
        rom[4][937] = 16'h0000;
        rom[4][938] = 16'h0000;
        rom[4][939] = 16'h0000;
        rom[4][940] = 16'h0000;
        rom[4][941] = 16'h0000;
        rom[4][942] = 16'h0000;
        rom[4][943] = 16'h0000;
        rom[4][944] = 16'h0000;
        rom[4][945] = 16'h0000;
        rom[4][946] = 16'h0000;
        rom[4][947] = 16'h0000;
        rom[4][948] = 16'h0000;
        rom[4][949] = 16'h0000;
        rom[4][950] = 16'h0000;
        rom[4][951] = 16'h0000;
        rom[4][952] = 16'h0000;
        rom[4][953] = 16'h0000;
        rom[4][954] = 16'h0000;
        rom[4][955] = 16'h0000;
        rom[4][956] = 16'h0000;
        rom[4][957] = 16'h0000;
        rom[4][958] = 16'h0000;
        rom[4][959] = 16'h0000;
        rom[4][960] = 16'h0000;
        rom[4][961] = 16'h0000;
        rom[4][962] = 16'h0000;
        rom[4][963] = 16'h0000;
        rom[4][964] = 16'h0000;
        rom[4][965] = 16'h0000;
        rom[4][966] = 16'h0000;
        rom[4][967] = 16'h0000;
        rom[4][968] = 16'h0000;
        rom[4][969] = 16'h0000;
        rom[4][970] = 16'h0000;
        rom[4][971] = 16'h0000;
        rom[4][972] = 16'h0000;
        rom[4][973] = 16'h0000;
        rom[4][974] = 16'h0000;
        rom[4][975] = 16'h0000;
        rom[4][976] = 16'h0000;
        rom[4][977] = 16'h0000;
        rom[4][978] = 16'h0000;
        rom[4][979] = 16'h0000;
        rom[4][980] = 16'hFF27;
        rom[4][981] = 16'hFE5D;
        rom[4][982] = 16'hFD7E;
        rom[4][983] = 16'hFE0E;
        rom[4][984] = 16'hFE6C;
        rom[4][985] = 16'hFE89;
        rom[4][986] = 16'hFEDF;
        rom[4][987] = 16'hFF3D;
        rom[4][988] = 16'h0024;
        rom[4][989] = 16'h01A3;
        rom[4][990] = 16'h0136;
        rom[4][991] = 16'h01A3;
        rom[4][992] = 16'h0169;
        rom[4][993] = 16'h00E7;
        rom[4][994] = 16'h00AD;
        rom[4][995] = 16'h0007;
        rom[4][996] = 16'hFFC6;
        rom[4][997] = 16'h0024;
        rom[4][998] = 16'hFF68;
        rom[4][999] = 16'hFF68;
        rom[4][1000] = 16'hFF19;
        rom[4][1001] = 16'hFECA;
        rom[4][1002] = 16'hFEDF;
        rom[4][1003] = 16'hFEBB;
        rom[4][1004] = 16'hFF20;
        rom[4][1005] = 16'hFEEE;
        rom[4][1006] = 16'hFF0B;
        rom[4][1007] = 16'hFEE7;
        rom[4][1008] = 16'hFED1;
        rom[4][1009] = 16'hFEF5;
        rom[4][1010] = 16'hFE65;
        rom[4][1011] = 16'hFDB0;
        rom[4][1012] = 16'h0000;
        rom[4][1013] = 16'h0000;
        rom[4][1014] = 16'h0000;
        rom[4][1015] = 16'h0000;
        rom[4][1016] = 16'h0000;
        rom[4][1017] = 16'h0000;
        rom[4][1018] = 16'h0000;
        rom[4][1019] = 16'h0000;
        rom[4][1020] = 16'h0000;
        rom[4][1021] = 16'h0000;
        rom[4][1022] = 16'h0000;
        rom[4][1023] = 16'h0000;
        rom[4][1024] = 16'h0000;
        rom[4][1025] = 16'h0000;
        rom[4][1026] = 16'h0000;
        rom[4][1027] = 16'h0000;
        rom[4][1028] = 16'h0000;
        rom[4][1029] = 16'h0000;
        rom[4][1030] = 16'h0000;
        rom[4][1031] = 16'h0000;
        rom[4][1032] = 16'h0000;
        rom[4][1033] = 16'h0000;
        rom[4][1034] = 16'h0000;
        rom[4][1035] = 16'h0000;
        rom[4][1036] = 16'h0000;
        rom[4][1037] = 16'h0000;
        rom[4][1038] = 16'h0000;
        rom[4][1039] = 16'h0000;
        rom[4][1040] = 16'h0000;
        rom[4][1041] = 16'h0000;
        rom[4][1042] = 16'h0000;
        rom[4][1043] = 16'h0000;
        rom[4][1044] = 16'h0000;
        rom[4][1045] = 16'h0000;
        rom[4][1046] = 16'h0000;
        rom[4][1047] = 16'h0000;
        rom[4][1048] = 16'h0000;
        rom[4][1049] = 16'h0000;
        rom[4][1050] = 16'h0000;
        rom[4][1051] = 16'h0000;
        rom[4][1052] = 16'h0000;
        rom[4][1053] = 16'h0000;
        rom[4][1054] = 16'h0000;
        rom[4][1055] = 16'h0000;
        rom[4][1056] = 16'h0000;
        rom[4][1057] = 16'h0000;
        rom[4][1058] = 16'h0000;
        rom[4][1059] = 16'h0000;
        rom[4][1060] = 16'h0000;
        rom[4][1061] = 16'h0000;
        rom[4][1062] = 16'h0000;
        rom[4][1063] = 16'h0000;
        rom[4][1064] = 16'h0000;
        rom[4][1065] = 16'h0000;
        rom[4][1066] = 16'h0000;
        rom[4][1067] = 16'h0000;
        rom[4][1068] = 16'h0000;
        rom[4][1069] = 16'h0000;
        rom[4][1070] = 16'h0000;
        rom[4][1071] = 16'h0000;
        rom[4][1072] = 16'h0000;
        rom[4][1073] = 16'h0000;
        rom[4][1074] = 16'h0000;
        rom[4][1075] = 16'h0000;
        rom[4][1076] = 16'h0000;
        rom[4][1077] = 16'h0000;
        rom[4][1078] = 16'hFFEA;
        rom[4][1079] = 16'hFF44;
        rom[4][1080] = 16'hFE56;
        rom[4][1081] = 16'hFF0B;
        rom[4][1082] = 16'hFFA9;
        rom[4][1083] = 16'h0007;
        rom[4][1084] = 16'h0016;
        rom[4][1085] = 16'h0033;
        rom[4][1086] = 16'h012F;
        rom[4][1087] = 16'h00D9;
        rom[4][1088] = 16'h00C3;
        rom[4][1089] = 16'h00E0;
        rom[4][1090] = 16'h00CA;
        rom[4][1091] = 16'h00B4;
        rom[4][1092] = 16'h00CA;
        rom[4][1093] = 16'h0136;
        rom[4][1094] = 16'h010B;
        rom[4][1095] = 16'h0098;
        rom[4][1096] = 16'hFFA9;
        rom[4][1097] = 16'h004F;
        rom[4][1098] = 16'h0098;
        rom[4][1099] = 16'h001D;
        rom[4][1100] = 16'hFF85;
        rom[4][1101] = 16'hFF27;
        rom[4][1102] = 16'hFF20;
        rom[4][1103] = 16'hFF44;
        rom[4][1104] = 16'hFF8D;
        rom[4][1105] = 16'hFF4C;
        rom[4][1106] = 16'hFF8D;
        rom[4][1107] = 16'h007B;
        rom[4][1108] = 16'hFFA9;
        rom[4][1109] = 16'hFF3D;
        rom[4][1110] = 16'h0000;
        rom[4][1111] = 16'h0000;
        rom[4][1112] = 16'h0000;
        rom[4][1113] = 16'h0000;
        rom[4][1114] = 16'h0000;
        rom[4][1115] = 16'h0000;
        rom[4][1116] = 16'h0000;
        rom[4][1117] = 16'h0000;
        rom[4][1118] = 16'h0000;
        rom[4][1119] = 16'h0000;
        rom[4][1120] = 16'h0000;
        rom[4][1121] = 16'h0000;
        rom[4][1122] = 16'h0000;
        rom[4][1123] = 16'h0000;
        rom[4][1124] = 16'h0000;
        rom[4][1125] = 16'h0000;
        rom[4][1126] = 16'h0000;
        rom[4][1127] = 16'h0000;
        rom[4][1128] = 16'h0000;
        rom[4][1129] = 16'h0000;
        rom[4][1130] = 16'h0000;
        rom[4][1131] = 16'h0000;
        rom[4][1132] = 16'h0000;
        rom[4][1133] = 16'h0000;
        rom[4][1134] = 16'h0000;
        rom[4][1135] = 16'h0000;
        rom[4][1136] = 16'h0000;
        rom[4][1137] = 16'h0000;
        rom[4][1138] = 16'h0000;
        rom[4][1139] = 16'h0000;
        rom[4][1140] = 16'h0000;
        rom[4][1141] = 16'h0000;
        rom[4][1142] = 16'h0000;
        rom[4][1143] = 16'h0000;
        rom[4][1144] = 16'h0000;
        rom[4][1145] = 16'h0000;
        rom[4][1146] = 16'h0000;
        rom[4][1147] = 16'h0000;
        rom[4][1148] = 16'h0000;
        rom[4][1149] = 16'h0000;
        rom[4][1150] = 16'h0000;
        rom[4][1151] = 16'h0000;
        rom[4][1152] = 16'h0000;
        rom[4][1153] = 16'h0000;
        rom[4][1154] = 16'h0000;
        rom[4][1155] = 16'h0000;
        rom[4][1156] = 16'h0000;
        rom[4][1157] = 16'h0000;
        rom[4][1158] = 16'h0000;
        rom[4][1159] = 16'h0000;
        rom[4][1160] = 16'h0000;
        rom[4][1161] = 16'h0000;
        rom[4][1162] = 16'h0000;
        rom[4][1163] = 16'h0000;
        rom[4][1164] = 16'h0000;
        rom[4][1165] = 16'h0000;
        rom[4][1166] = 16'h0000;
        rom[4][1167] = 16'h0000;
        rom[4][1168] = 16'h0000;
        rom[4][1169] = 16'h0000;
        rom[4][1170] = 16'h0000;
        rom[4][1171] = 16'h0000;
        rom[4][1172] = 16'h0000;
        rom[4][1173] = 16'h0000;
        rom[4][1174] = 16'h0000;
        rom[4][1175] = 16'h0000;
        rom[4][1176] = 16'hFF7E;
        rom[4][1177] = 16'hFEE7;
        rom[4][1178] = 16'hFE32;
        rom[4][1179] = 16'hFE97;
        rom[4][1180] = 16'hFFA9;
        rom[4][1181] = 16'h0000;
        rom[4][1182] = 16'hFFC6;
        rom[4][1183] = 16'hFF85;
        rom[4][1184] = 16'hFF20;
        rom[4][1185] = 16'hFEF5;
        rom[4][1186] = 16'hFEA6;
        rom[4][1187] = 16'hFE24;
        rom[4][1188] = 16'hFDE3;
        rom[4][1189] = 16'hFE0E;
        rom[4][1190] = 16'hFED1;
        rom[4][1191] = 16'hFFA2;
        rom[4][1192] = 16'hFFB1;
        rom[4][1193] = 16'hFF94;
        rom[4][1194] = 16'hFF9B;
        rom[4][1195] = 16'hFF8D;
        rom[4][1196] = 16'hFF9B;
        rom[4][1197] = 16'hFF77;
        rom[4][1198] = 16'hFF20;
        rom[4][1199] = 16'hFF4C;
        rom[4][1200] = 16'hFF70;
        rom[4][1201] = 16'hFF44;
        rom[4][1202] = 16'hFF8D;
        rom[4][1203] = 16'hFF36;
        rom[4][1204] = 16'hFF5A;
        rom[4][1205] = 16'hFF70;
        rom[4][1206] = 16'hFEFC;
        rom[4][1207] = 16'hFF4C;
        rom[4][1208] = 16'h0000;
        rom[4][1209] = 16'h0000;
        rom[4][1210] = 16'h0000;
        rom[4][1211] = 16'h0000;
        rom[4][1212] = 16'h0000;
        rom[4][1213] = 16'h0000;
        rom[4][1214] = 16'h0000;
        rom[4][1215] = 16'h0000;
        rom[4][1216] = 16'h0000;
        rom[4][1217] = 16'h0000;
        rom[4][1218] = 16'h0000;
        rom[4][1219] = 16'h0000;
        rom[4][1220] = 16'h0000;
        rom[4][1221] = 16'h0000;
        rom[4][1222] = 16'h0000;
        rom[4][1223] = 16'h0000;
        rom[4][1224] = 16'h0000;
        rom[4][1225] = 16'h0000;
        rom[4][1226] = 16'h0000;
        rom[4][1227] = 16'h0000;
        rom[4][1228] = 16'h0000;
        rom[4][1229] = 16'h0000;
        rom[4][1230] = 16'h0000;
        rom[4][1231] = 16'h0000;
        rom[4][1232] = 16'h0000;
        rom[4][1233] = 16'h0000;
        rom[4][1234] = 16'h0000;
        rom[4][1235] = 16'h0000;
        rom[4][1236] = 16'h0000;
        rom[4][1237] = 16'h0000;
        rom[4][1238] = 16'h0000;
        rom[4][1239] = 16'h0000;
        rom[4][1240] = 16'h0000;
        rom[4][1241] = 16'h0000;
        rom[4][1242] = 16'h0000;
        rom[4][1243] = 16'h0000;
        rom[4][1244] = 16'h0000;
        rom[4][1245] = 16'h0000;
        rom[4][1246] = 16'h0000;
        rom[4][1247] = 16'h0000;
        rom[4][1248] = 16'h0000;
        rom[4][1249] = 16'h0000;
        rom[4][1250] = 16'h0000;
        rom[4][1251] = 16'h0000;
        rom[4][1252] = 16'h0000;
        rom[4][1253] = 16'h0000;
        rom[4][1254] = 16'h0000;
        rom[4][1255] = 16'h0000;
        rom[4][1256] = 16'h0000;
        rom[4][1257] = 16'h0000;
        rom[4][1258] = 16'h0000;
        rom[4][1259] = 16'h0000;
        rom[4][1260] = 16'h0000;
        rom[4][1261] = 16'h0000;
        rom[4][1262] = 16'h0000;
        rom[4][1263] = 16'h0000;
        rom[4][1264] = 16'h0000;
        rom[4][1265] = 16'h0000;
        rom[4][1266] = 16'h0000;
        rom[4][1267] = 16'h0000;
        rom[4][1268] = 16'h0000;
        rom[4][1269] = 16'h0000;
        rom[4][1270] = 16'h0000;
        rom[4][1271] = 16'h0000;
        rom[4][1272] = 16'h0000;
        rom[4][1273] = 16'h0000;
        rom[5][0] = 16'hFFA9;
        rom[5][1] = 16'hFFA9;
        rom[5][2] = 16'hFF9B;
        rom[5][3] = 16'hFF94;
        rom[5][4] = 16'h0024;
        rom[5][5] = 16'h00AD;
        rom[5][6] = 16'h00E7;
        rom[5][7] = 16'h012F;
        rom[5][8] = 16'h0136;
        rom[5][9] = 16'h0112;
        rom[5][10] = 16'h00EE;
        rom[5][11] = 16'h00CA;
        rom[5][12] = 16'h00B4;
        rom[5][13] = 16'h009F;
        rom[5][14] = 16'h0082;
        rom[5][15] = 16'h007B;
        rom[5][16] = 16'h005E;
        rom[5][17] = 16'h0024;
        rom[5][18] = 16'hFFE3;
        rom[5][19] = 16'hFFA2;
        rom[5][20] = 16'hFF7E;
        rom[5][21] = 16'hFF61;
        rom[5][22] = 16'hFF3D;
        rom[5][23] = 16'hFF36;
        rom[5][24] = 16'hFF3D;
        rom[5][25] = 16'hFF53;
        rom[5][26] = 16'hFF68;
        rom[5][27] = 16'hFF77;
        rom[5][28] = 16'hFF94;
        rom[5][29] = 16'hFFA9;
        rom[5][30] = 16'hFFBF;
        rom[5][31] = 16'hFFC6;
        rom[5][32] = 16'h0000;
        rom[5][33] = 16'h0000;
        rom[5][34] = 16'h0000;
        rom[5][35] = 16'h0000;
        rom[5][36] = 16'h0000;
        rom[5][37] = 16'h0000;
        rom[5][38] = 16'h0000;
        rom[5][39] = 16'h0000;
        rom[5][40] = 16'h0000;
        rom[5][41] = 16'h0000;
        rom[5][42] = 16'h0000;
        rom[5][43] = 16'h0000;
        rom[5][44] = 16'h0000;
        rom[5][45] = 16'h0000;
        rom[5][46] = 16'h0000;
        rom[5][47] = 16'h0000;
        rom[5][48] = 16'h0000;
        rom[5][49] = 16'h0000;
        rom[5][50] = 16'h0000;
        rom[5][51] = 16'h0000;
        rom[5][52] = 16'h0000;
        rom[5][53] = 16'h0000;
        rom[5][54] = 16'h0000;
        rom[5][55] = 16'h0000;
        rom[5][56] = 16'h0000;
        rom[5][57] = 16'h0000;
        rom[5][58] = 16'h0000;
        rom[5][59] = 16'h0000;
        rom[5][60] = 16'h0000;
        rom[5][61] = 16'h0000;
        rom[5][62] = 16'h0000;
        rom[5][63] = 16'h0000;
        rom[5][64] = 16'h0000;
        rom[5][65] = 16'h0000;
        rom[5][66] = 16'h0000;
        rom[5][67] = 16'h0000;
        rom[5][68] = 16'h0000;
        rom[5][69] = 16'h0000;
        rom[5][70] = 16'h0000;
        rom[5][71] = 16'h0000;
        rom[5][72] = 16'h0000;
        rom[5][73] = 16'h0000;
        rom[5][74] = 16'h0000;
        rom[5][75] = 16'h0000;
        rom[5][76] = 16'h0000;
        rom[5][77] = 16'h0000;
        rom[5][78] = 16'h0000;
        rom[5][79] = 16'h0000;
        rom[5][80] = 16'h0000;
        rom[5][81] = 16'h0000;
        rom[5][82] = 16'h0000;
        rom[5][83] = 16'h0000;
        rom[5][84] = 16'h0000;
        rom[5][85] = 16'h0000;
        rom[5][86] = 16'h0000;
        rom[5][87] = 16'h0000;
        rom[5][88] = 16'h0000;
        rom[5][89] = 16'h0000;
        rom[5][90] = 16'h0000;
        rom[5][91] = 16'h0000;
        rom[5][92] = 16'h0000;
        rom[5][93] = 16'h0000;
        rom[5][94] = 16'h0000;
        rom[5][95] = 16'h0000;
        rom[5][96] = 16'h0000;
        rom[5][97] = 16'h0000;
        rom[5][98] = 16'h00AD;
        rom[5][99] = 16'h00CA;
        rom[5][100] = 16'h009F;
        rom[5][101] = 16'h0098;
        rom[5][102] = 16'h013E;
        rom[5][103] = 16'h010B;
        rom[5][104] = 16'h00CA;
        rom[5][105] = 16'h00D1;
        rom[5][106] = 16'h00BC;
        rom[5][107] = 16'h009F;
        rom[5][108] = 16'h0090;
        rom[5][109] = 16'h0098;
        rom[5][110] = 16'h0089;
        rom[5][111] = 16'h0090;
        rom[5][112] = 16'h00A6;
        rom[5][113] = 16'h00AD;
        rom[5][114] = 16'h00BC;
        rom[5][115] = 16'h00E0;
        rom[5][116] = 16'h00E7;
        rom[5][117] = 16'h00D1;
        rom[5][118] = 16'h009F;
        rom[5][119] = 16'h0089;
        rom[5][120] = 16'h003A;
        rom[5][121] = 16'h000E;
        rom[5][122] = 16'h001D;
        rom[5][123] = 16'h002B;
        rom[5][124] = 16'h0033;
        rom[5][125] = 16'h0048;
        rom[5][126] = 16'h007B;
        rom[5][127] = 16'h009F;
        rom[5][128] = 16'h00A6;
        rom[5][129] = 16'h00AD;
        rom[5][130] = 16'h0000;
        rom[5][131] = 16'h0000;
        rom[5][132] = 16'h0000;
        rom[5][133] = 16'h0000;
        rom[5][134] = 16'h0000;
        rom[5][135] = 16'h0000;
        rom[5][136] = 16'h0000;
        rom[5][137] = 16'h0000;
        rom[5][138] = 16'h0000;
        rom[5][139] = 16'h0000;
        rom[5][140] = 16'h0000;
        rom[5][141] = 16'h0000;
        rom[5][142] = 16'h0000;
        rom[5][143] = 16'h0000;
        rom[5][144] = 16'h0000;
        rom[5][145] = 16'h0000;
        rom[5][146] = 16'h0000;
        rom[5][147] = 16'h0000;
        rom[5][148] = 16'h0000;
        rom[5][149] = 16'h0000;
        rom[5][150] = 16'h0000;
        rom[5][151] = 16'h0000;
        rom[5][152] = 16'h0000;
        rom[5][153] = 16'h0000;
        rom[5][154] = 16'h0000;
        rom[5][155] = 16'h0000;
        rom[5][156] = 16'h0000;
        rom[5][157] = 16'h0000;
        rom[5][158] = 16'h0000;
        rom[5][159] = 16'h0000;
        rom[5][160] = 16'h0000;
        rom[5][161] = 16'h0000;
        rom[5][162] = 16'h0000;
        rom[5][163] = 16'h0000;
        rom[5][164] = 16'h0000;
        rom[5][165] = 16'h0000;
        rom[5][166] = 16'h0000;
        rom[5][167] = 16'h0000;
        rom[5][168] = 16'h0000;
        rom[5][169] = 16'h0000;
        rom[5][170] = 16'h0000;
        rom[5][171] = 16'h0000;
        rom[5][172] = 16'h0000;
        rom[5][173] = 16'h0000;
        rom[5][174] = 16'h0000;
        rom[5][175] = 16'h0000;
        rom[5][176] = 16'h0000;
        rom[5][177] = 16'h0000;
        rom[5][178] = 16'h0000;
        rom[5][179] = 16'h0000;
        rom[5][180] = 16'h0000;
        rom[5][181] = 16'h0000;
        rom[5][182] = 16'h0000;
        rom[5][183] = 16'h0000;
        rom[5][184] = 16'h0000;
        rom[5][185] = 16'h0000;
        rom[5][186] = 16'h0000;
        rom[5][187] = 16'h0000;
        rom[5][188] = 16'h0000;
        rom[5][189] = 16'h0000;
        rom[5][190] = 16'h0000;
        rom[5][191] = 16'h0000;
        rom[5][192] = 16'h0000;
        rom[5][193] = 16'h0000;
        rom[5][194] = 16'h0000;
        rom[5][195] = 16'h0000;
        rom[5][196] = 16'h003A;
        rom[5][197] = 16'h0024;
        rom[5][198] = 16'h0024;
        rom[5][199] = 16'h0041;
        rom[5][200] = 16'h00FD;
        rom[5][201] = 16'h005E;
        rom[5][202] = 16'hFFE3;
        rom[5][203] = 16'hFF7E;
        rom[5][204] = 16'hFF5A;
        rom[5][205] = 16'hFF3D;
        rom[5][206] = 16'hFF4C;
        rom[5][207] = 16'hFF36;
        rom[5][208] = 16'hFF27;
        rom[5][209] = 16'hFF61;
        rom[5][210] = 16'hFFA2;
        rom[5][211] = 16'hFFCD;
        rom[5][212] = 16'hFFF9;
        rom[5][213] = 16'h0041;
        rom[5][214] = 16'h009F;
        rom[5][215] = 16'h00FD;
        rom[5][216] = 16'h00E0;
        rom[5][217] = 16'h0089;
        rom[5][218] = 16'h0057;
        rom[5][219] = 16'h0048;
        rom[5][220] = 16'h0048;
        rom[5][221] = 16'h003A;
        rom[5][222] = 16'h000E;
        rom[5][223] = 16'h001D;
        rom[5][224] = 16'h004F;
        rom[5][225] = 16'h0048;
        rom[5][226] = 16'h0007;
        rom[5][227] = 16'h002B;
        rom[5][228] = 16'h0000;
        rom[5][229] = 16'h0000;
        rom[5][230] = 16'h0000;
        rom[5][231] = 16'h0000;
        rom[5][232] = 16'h0000;
        rom[5][233] = 16'h0000;
        rom[5][234] = 16'h0000;
        rom[5][235] = 16'h0000;
        rom[5][236] = 16'h0000;
        rom[5][237] = 16'h0000;
        rom[5][238] = 16'h0000;
        rom[5][239] = 16'h0000;
        rom[5][240] = 16'h0000;
        rom[5][241] = 16'h0000;
        rom[5][242] = 16'h0000;
        rom[5][243] = 16'h0000;
        rom[5][244] = 16'h0000;
        rom[5][245] = 16'h0000;
        rom[5][246] = 16'h0000;
        rom[5][247] = 16'h0000;
        rom[5][248] = 16'h0000;
        rom[5][249] = 16'h0000;
        rom[5][250] = 16'h0000;
        rom[5][251] = 16'h0000;
        rom[5][252] = 16'h0000;
        rom[5][253] = 16'h0000;
        rom[5][254] = 16'h0000;
        rom[5][255] = 16'h0000;
        rom[5][256] = 16'h0000;
        rom[5][257] = 16'h0000;
        rom[5][258] = 16'h0000;
        rom[5][259] = 16'h0000;
        rom[5][260] = 16'h0000;
        rom[5][261] = 16'h0000;
        rom[5][262] = 16'h0000;
        rom[5][263] = 16'h0000;
        rom[5][264] = 16'h0000;
        rom[5][265] = 16'h0000;
        rom[5][266] = 16'h0000;
        rom[5][267] = 16'h0000;
        rom[5][268] = 16'h0000;
        rom[5][269] = 16'h0000;
        rom[5][270] = 16'h0000;
        rom[5][271] = 16'h0000;
        rom[5][272] = 16'h0000;
        rom[5][273] = 16'h0000;
        rom[5][274] = 16'h0000;
        rom[5][275] = 16'h0000;
        rom[5][276] = 16'h0000;
        rom[5][277] = 16'h0000;
        rom[5][278] = 16'h0000;
        rom[5][279] = 16'h0000;
        rom[5][280] = 16'h0000;
        rom[5][281] = 16'h0000;
        rom[5][282] = 16'h0000;
        rom[5][283] = 16'h0000;
        rom[5][284] = 16'h0000;
        rom[5][285] = 16'h0000;
        rom[5][286] = 16'h0000;
        rom[5][287] = 16'h0000;
        rom[5][288] = 16'h0000;
        rom[5][289] = 16'h0000;
        rom[5][290] = 16'h0000;
        rom[5][291] = 16'h0000;
        rom[5][292] = 16'h0000;
        rom[5][293] = 16'h0000;
        rom[5][294] = 16'hFEBB;
        rom[5][295] = 16'hFF03;
        rom[5][296] = 16'hFF70;
        rom[5][297] = 16'hFFB1;
        rom[5][298] = 16'h0162;
        rom[5][299] = 16'h02CB;
        rom[5][300] = 16'h02E7;
        rom[5][301] = 16'h01C7;
        rom[5][302] = 16'h00FD;
        rom[5][303] = 16'h0073;
        rom[5][304] = 16'h003A;
        rom[5][305] = 16'h002B;
        rom[5][306] = 16'h005E;
        rom[5][307] = 16'h005E;
        rom[5][308] = 16'h004F;
        rom[5][309] = 16'h006C;
        rom[5][310] = 16'h005E;
        rom[5][311] = 16'h0065;
        rom[5][312] = 16'h0098;
        rom[5][313] = 16'h00AD;
        rom[5][314] = 16'h006C;
        rom[5][315] = 16'hFFF9;
        rom[5][316] = 16'hFFF2;
        rom[5][317] = 16'h0024;
        rom[5][318] = 16'hFFF9;
        rom[5][319] = 16'hFFF9;
        rom[5][320] = 16'hFFEA;
        rom[5][321] = 16'hFFCD;
        rom[5][322] = 16'hFFC6;
        rom[5][323] = 16'hFF77;
        rom[5][324] = 16'hFF53;
        rom[5][325] = 16'hFF3D;
        rom[5][326] = 16'h0000;
        rom[5][327] = 16'h0000;
        rom[5][328] = 16'h0000;
        rom[5][329] = 16'h0000;
        rom[5][330] = 16'h0000;
        rom[5][331] = 16'h0000;
        rom[5][332] = 16'h0000;
        rom[5][333] = 16'h0000;
        rom[5][334] = 16'h0000;
        rom[5][335] = 16'h0000;
        rom[5][336] = 16'h0000;
        rom[5][337] = 16'h0000;
        rom[5][338] = 16'h0000;
        rom[5][339] = 16'h0000;
        rom[5][340] = 16'h0000;
        rom[5][341] = 16'h0000;
        rom[5][342] = 16'h0000;
        rom[5][343] = 16'h0000;
        rom[5][344] = 16'h0000;
        rom[5][345] = 16'h0000;
        rom[5][346] = 16'h0000;
        rom[5][347] = 16'h0000;
        rom[5][348] = 16'h0000;
        rom[5][349] = 16'h0000;
        rom[5][350] = 16'h0000;
        rom[5][351] = 16'h0000;
        rom[5][352] = 16'h0000;
        rom[5][353] = 16'h0000;
        rom[5][354] = 16'h0000;
        rom[5][355] = 16'h0000;
        rom[5][356] = 16'h0000;
        rom[5][357] = 16'h0000;
        rom[5][358] = 16'h0000;
        rom[5][359] = 16'h0000;
        rom[5][360] = 16'h0000;
        rom[5][361] = 16'h0000;
        rom[5][362] = 16'h0000;
        rom[5][363] = 16'h0000;
        rom[5][364] = 16'h0000;
        rom[5][365] = 16'h0000;
        rom[5][366] = 16'h0000;
        rom[5][367] = 16'h0000;
        rom[5][368] = 16'h0000;
        rom[5][369] = 16'h0000;
        rom[5][370] = 16'h0000;
        rom[5][371] = 16'h0000;
        rom[5][372] = 16'h0000;
        rom[5][373] = 16'h0000;
        rom[5][374] = 16'h0000;
        rom[5][375] = 16'h0000;
        rom[5][376] = 16'h0000;
        rom[5][377] = 16'h0000;
        rom[5][378] = 16'h0000;
        rom[5][379] = 16'h0000;
        rom[5][380] = 16'h0000;
        rom[5][381] = 16'h0000;
        rom[5][382] = 16'h0000;
        rom[5][383] = 16'h0000;
        rom[5][384] = 16'h0000;
        rom[5][385] = 16'h0000;
        rom[5][386] = 16'h0000;
        rom[5][387] = 16'h0000;
        rom[5][388] = 16'h0000;
        rom[5][389] = 16'h0000;
        rom[5][390] = 16'h0000;
        rom[5][391] = 16'h0000;
        rom[5][392] = 16'hFEFC;
        rom[5][393] = 16'hFF70;
        rom[5][394] = 16'h0000;
        rom[5][395] = 16'h0033;
        rom[5][396] = 16'h00D1;
        rom[5][397] = 16'h005E;
        rom[5][398] = 16'hFFB8;
        rom[5][399] = 16'hFE73;
        rom[5][400] = 16'hFE56;
        rom[5][401] = 16'hFE65;
        rom[5][402] = 16'hFE5D;
        rom[5][403] = 16'hFE4F;
        rom[5][404] = 16'hFE6C;
        rom[5][405] = 16'hFE56;
        rom[5][406] = 16'hFE5D;
        rom[5][407] = 16'hFE81;
        rom[5][408] = 16'hFEB4;
        rom[5][409] = 16'hFED1;
        rom[5][410] = 16'hFEEE;
        rom[5][411] = 16'hFF27;
        rom[5][412] = 16'hFFA2;
        rom[5][413] = 16'h0000;
        rom[5][414] = 16'h001D;
        rom[5][415] = 16'h0065;
        rom[5][416] = 16'h0057;
        rom[5][417] = 16'h0065;
        rom[5][418] = 16'h005E;
        rom[5][419] = 16'hFFF9;
        rom[5][420] = 16'h0007;
        rom[5][421] = 16'hFFB8;
        rom[5][422] = 16'hFF70;
        rom[5][423] = 16'hFF4C;
        rom[5][424] = 16'h0000;
        rom[5][425] = 16'h0000;
        rom[5][426] = 16'h0000;
        rom[5][427] = 16'h0000;
        rom[5][428] = 16'h0000;
        rom[5][429] = 16'h0000;
        rom[5][430] = 16'h0000;
        rom[5][431] = 16'h0000;
        rom[5][432] = 16'h0000;
        rom[5][433] = 16'h0000;
        rom[5][434] = 16'h0000;
        rom[5][435] = 16'h0000;
        rom[5][436] = 16'h0000;
        rom[5][437] = 16'h0000;
        rom[5][438] = 16'h0000;
        rom[5][439] = 16'h0000;
        rom[5][440] = 16'h0000;
        rom[5][441] = 16'h0000;
        rom[5][442] = 16'h0000;
        rom[5][443] = 16'h0000;
        rom[5][444] = 16'h0000;
        rom[5][445] = 16'h0000;
        rom[5][446] = 16'h0000;
        rom[5][447] = 16'h0000;
        rom[5][448] = 16'h0000;
        rom[5][449] = 16'h0000;
        rom[5][450] = 16'h0000;
        rom[5][451] = 16'h0000;
        rom[5][452] = 16'h0000;
        rom[5][453] = 16'h0000;
        rom[5][454] = 16'h0000;
        rom[5][455] = 16'h0000;
        rom[5][456] = 16'h0000;
        rom[5][457] = 16'h0000;
        rom[5][458] = 16'h0000;
        rom[5][459] = 16'h0000;
        rom[5][460] = 16'h0000;
        rom[5][461] = 16'h0000;
        rom[5][462] = 16'h0000;
        rom[5][463] = 16'h0000;
        rom[5][464] = 16'h0000;
        rom[5][465] = 16'h0000;
        rom[5][466] = 16'h0000;
        rom[5][467] = 16'h0000;
        rom[5][468] = 16'h0000;
        rom[5][469] = 16'h0000;
        rom[5][470] = 16'h0000;
        rom[5][471] = 16'h0000;
        rom[5][472] = 16'h0000;
        rom[5][473] = 16'h0000;
        rom[5][474] = 16'h0000;
        rom[5][475] = 16'h0000;
        rom[5][476] = 16'h0000;
        rom[5][477] = 16'h0000;
        rom[5][478] = 16'h0000;
        rom[5][479] = 16'h0000;
        rom[5][480] = 16'h0000;
        rom[5][481] = 16'h0000;
        rom[5][482] = 16'h0000;
        rom[5][483] = 16'h0000;
        rom[5][484] = 16'h0000;
        rom[5][485] = 16'h0000;
        rom[5][486] = 16'h0000;
        rom[5][487] = 16'h0000;
        rom[5][488] = 16'h0000;
        rom[5][489] = 16'h0000;
        rom[5][490] = 16'hFFB8;
        rom[5][491] = 16'hFFD5;
        rom[5][492] = 16'h001D;
        rom[5][493] = 16'h001D;
        rom[5][494] = 16'h000E;
        rom[5][495] = 16'h0057;
        rom[5][496] = 16'h00F5;
        rom[5][497] = 16'h014C;
        rom[5][498] = 16'h019B;
        rom[5][499] = 16'h01CE;
        rom[5][500] = 16'h01B1;
        rom[5][501] = 16'h0194;
        rom[5][502] = 16'h01B8;
        rom[5][503] = 16'h01AA;
        rom[5][504] = 16'h017F;
        rom[5][505] = 16'h0177;
        rom[5][506] = 16'h018D;
        rom[5][507] = 16'h0145;
        rom[5][508] = 16'h00CA;
        rom[5][509] = 16'h00EE;
        rom[5][510] = 16'h0112;
        rom[5][511] = 16'h00E7;
        rom[5][512] = 16'h0073;
        rom[5][513] = 16'h0090;
        rom[5][514] = 16'h003A;
        rom[5][515] = 16'hFFF9;
        rom[5][516] = 16'h000E;
        rom[5][517] = 16'h0016;
        rom[5][518] = 16'h0041;
        rom[5][519] = 16'h0016;
        rom[5][520] = 16'hFFE3;
        rom[5][521] = 16'hFFEA;
        rom[5][522] = 16'h0000;
        rom[5][523] = 16'h0000;
        rom[5][524] = 16'h0000;
        rom[5][525] = 16'h0000;
        rom[5][526] = 16'h0000;
        rom[5][527] = 16'h0000;
        rom[5][528] = 16'h0000;
        rom[5][529] = 16'h0000;
        rom[5][530] = 16'h0000;
        rom[5][531] = 16'h0000;
        rom[5][532] = 16'h0000;
        rom[5][533] = 16'h0000;
        rom[5][534] = 16'h0000;
        rom[5][535] = 16'h0000;
        rom[5][536] = 16'h0000;
        rom[5][537] = 16'h0000;
        rom[5][538] = 16'h0000;
        rom[5][539] = 16'h0000;
        rom[5][540] = 16'h0000;
        rom[5][541] = 16'h0000;
        rom[5][542] = 16'h0000;
        rom[5][543] = 16'h0000;
        rom[5][544] = 16'h0000;
        rom[5][545] = 16'h0000;
        rom[5][546] = 16'h0000;
        rom[5][547] = 16'h0000;
        rom[5][548] = 16'h0000;
        rom[5][549] = 16'h0000;
        rom[5][550] = 16'h0000;
        rom[5][551] = 16'h0000;
        rom[5][552] = 16'h0000;
        rom[5][553] = 16'h0000;
        rom[5][554] = 16'h0000;
        rom[5][555] = 16'h0000;
        rom[5][556] = 16'h0000;
        rom[5][557] = 16'h0000;
        rom[5][558] = 16'h0000;
        rom[5][559] = 16'h0000;
        rom[5][560] = 16'h0000;
        rom[5][561] = 16'h0000;
        rom[5][562] = 16'h0000;
        rom[5][563] = 16'h0000;
        rom[5][564] = 16'h0000;
        rom[5][565] = 16'h0000;
        rom[5][566] = 16'h0000;
        rom[5][567] = 16'h0000;
        rom[5][568] = 16'h0000;
        rom[5][569] = 16'h0000;
        rom[5][570] = 16'h0000;
        rom[5][571] = 16'h0000;
        rom[5][572] = 16'h0000;
        rom[5][573] = 16'h0000;
        rom[5][574] = 16'h0000;
        rom[5][575] = 16'h0000;
        rom[5][576] = 16'h0000;
        rom[5][577] = 16'h0000;
        rom[5][578] = 16'h0000;
        rom[5][579] = 16'h0000;
        rom[5][580] = 16'h0000;
        rom[5][581] = 16'h0000;
        rom[5][582] = 16'h0000;
        rom[5][583] = 16'h0000;
        rom[5][584] = 16'h0000;
        rom[5][585] = 16'h0000;
        rom[5][586] = 16'h0000;
        rom[5][587] = 16'h0000;
        rom[5][588] = 16'h0145;
        rom[5][589] = 16'h010B;
        rom[5][590] = 16'h00E7;
        rom[5][591] = 16'h00D1;
        rom[5][592] = 16'hFD7E;
        rom[5][593] = 16'h02FD;
        rom[5][594] = 16'h02D9;
        rom[5][595] = 16'h038D;
        rom[5][596] = 16'hFD2E;
        rom[5][597] = 16'hFE2B;
        rom[5][598] = 16'hFE65;
        rom[5][599] = 16'hFEA6;
        rom[5][600] = 16'hFEDF;
        rom[5][601] = 16'hFEE7;
        rom[5][602] = 16'hFEAD;
        rom[5][603] = 16'hFE41;
        rom[5][604] = 16'hFE73;
        rom[5][605] = 16'hFF0B;
        rom[5][606] = 16'hFFB1;
        rom[5][607] = 16'h006C;
        rom[5][608] = 16'h005E;
        rom[5][609] = 16'h005E;
        rom[5][610] = 16'h00BC;
        rom[5][611] = 16'h00E7;
        rom[5][612] = 16'h00E0;
        rom[5][613] = 16'h0112;
        rom[5][614] = 16'h0186;
        rom[5][615] = 16'h018D;
        rom[5][616] = 16'h0169;
        rom[5][617] = 16'h0194;
        rom[5][618] = 16'h0177;
        rom[5][619] = 16'h0145;
        rom[5][620] = 16'h0000;
        rom[5][621] = 16'h0000;
        rom[5][622] = 16'h0000;
        rom[5][623] = 16'h0000;
        rom[5][624] = 16'h0000;
        rom[5][625] = 16'h0000;
        rom[5][626] = 16'h0000;
        rom[5][627] = 16'h0000;
        rom[5][628] = 16'h0000;
        rom[5][629] = 16'h0000;
        rom[5][630] = 16'h0000;
        rom[5][631] = 16'h0000;
        rom[5][632] = 16'h0000;
        rom[5][633] = 16'h0000;
        rom[5][634] = 16'h0000;
        rom[5][635] = 16'h0000;
        rom[5][636] = 16'h0000;
        rom[5][637] = 16'h0000;
        rom[5][638] = 16'h0000;
        rom[5][639] = 16'h0000;
        rom[5][640] = 16'h0000;
        rom[5][641] = 16'h0000;
        rom[5][642] = 16'h0000;
        rom[5][643] = 16'h0000;
        rom[5][644] = 16'h0000;
        rom[5][645] = 16'h0000;
        rom[5][646] = 16'h0000;
        rom[5][647] = 16'h0000;
        rom[5][648] = 16'h0000;
        rom[5][649] = 16'h0000;
        rom[5][650] = 16'h0000;
        rom[5][651] = 16'h0000;
        rom[5][652] = 16'h0000;
        rom[5][653] = 16'h0000;
        rom[5][654] = 16'h0000;
        rom[5][655] = 16'h0000;
        rom[5][656] = 16'h0000;
        rom[5][657] = 16'h0000;
        rom[5][658] = 16'h0000;
        rom[5][659] = 16'h0000;
        rom[5][660] = 16'h0000;
        rom[5][661] = 16'h0000;
        rom[5][662] = 16'h0000;
        rom[5][663] = 16'h0000;
        rom[5][664] = 16'h0000;
        rom[5][665] = 16'h0000;
        rom[5][666] = 16'h0000;
        rom[5][667] = 16'h0000;
        rom[5][668] = 16'h0000;
        rom[5][669] = 16'h0000;
        rom[5][670] = 16'h0000;
        rom[5][671] = 16'h0000;
        rom[5][672] = 16'h0000;
        rom[5][673] = 16'h0000;
        rom[5][674] = 16'h0000;
        rom[5][675] = 16'h0000;
        rom[5][676] = 16'h0000;
        rom[5][677] = 16'h0000;
        rom[5][678] = 16'h0000;
        rom[5][679] = 16'h0000;
        rom[5][680] = 16'h0000;
        rom[5][681] = 16'h0000;
        rom[5][682] = 16'h0000;
        rom[5][683] = 16'h0000;
        rom[5][684] = 16'h0000;
        rom[5][685] = 16'h0000;
        rom[5][686] = 16'h0128;
        rom[5][687] = 16'h00AD;
        rom[5][688] = 16'h0048;
        rom[5][689] = 16'h004F;
        rom[5][690] = 16'hFFB1;
        rom[5][691] = 16'hFF9B;
        rom[5][692] = 16'hFF77;
        rom[5][693] = 16'hFF4C;
        rom[5][694] = 16'hFF12;
        rom[5][695] = 16'hFF44;
        rom[5][696] = 16'hFF85;
        rom[5][697] = 16'hFFB1;
        rom[5][698] = 16'hFFF9;
        rom[5][699] = 16'h0016;
        rom[5][700] = 16'h0041;
        rom[5][701] = 16'h0098;
        rom[5][702] = 16'h007B;
        rom[5][703] = 16'h007B;
        rom[5][704] = 16'h0065;
        rom[5][705] = 16'h006C;
        rom[5][706] = 16'h009F;
        rom[5][707] = 16'h0098;
        rom[5][708] = 16'h0082;
        rom[5][709] = 16'h006C;
        rom[5][710] = 16'h00E7;
        rom[5][711] = 16'h0112;
        rom[5][712] = 16'h0119;
        rom[5][713] = 16'h010B;
        rom[5][714] = 16'h010B;
        rom[5][715] = 16'h0153;
        rom[5][716] = 16'h0128;
        rom[5][717] = 16'h0098;
        rom[5][718] = 16'h0000;
        rom[5][719] = 16'h0000;
        rom[5][720] = 16'h0000;
        rom[5][721] = 16'h0000;
        rom[5][722] = 16'h0000;
        rom[5][723] = 16'h0000;
        rom[5][724] = 16'h0000;
        rom[5][725] = 16'h0000;
        rom[5][726] = 16'h0000;
        rom[5][727] = 16'h0000;
        rom[5][728] = 16'h0000;
        rom[5][729] = 16'h0000;
        rom[5][730] = 16'h0000;
        rom[5][731] = 16'h0000;
        rom[5][732] = 16'h0000;
        rom[5][733] = 16'h0000;
        rom[5][734] = 16'h0000;
        rom[5][735] = 16'h0000;
        rom[5][736] = 16'h0000;
        rom[5][737] = 16'h0000;
        rom[5][738] = 16'h0000;
        rom[5][739] = 16'h0000;
        rom[5][740] = 16'h0000;
        rom[5][741] = 16'h0000;
        rom[5][742] = 16'h0000;
        rom[5][743] = 16'h0000;
        rom[5][744] = 16'h0000;
        rom[5][745] = 16'h0000;
        rom[5][746] = 16'h0000;
        rom[5][747] = 16'h0000;
        rom[5][748] = 16'h0000;
        rom[5][749] = 16'h0000;
        rom[5][750] = 16'h0000;
        rom[5][751] = 16'h0000;
        rom[5][752] = 16'h0000;
        rom[5][753] = 16'h0000;
        rom[5][754] = 16'h0000;
        rom[5][755] = 16'h0000;
        rom[5][756] = 16'h0000;
        rom[5][757] = 16'h0000;
        rom[5][758] = 16'h0000;
        rom[5][759] = 16'h0000;
        rom[5][760] = 16'h0000;
        rom[5][761] = 16'h0000;
        rom[5][762] = 16'h0000;
        rom[5][763] = 16'h0000;
        rom[5][764] = 16'h0000;
        rom[5][765] = 16'h0000;
        rom[5][766] = 16'h0000;
        rom[5][767] = 16'h0000;
        rom[5][768] = 16'h0000;
        rom[5][769] = 16'h0000;
        rom[5][770] = 16'h0000;
        rom[5][771] = 16'h0000;
        rom[5][772] = 16'h0000;
        rom[5][773] = 16'h0000;
        rom[5][774] = 16'h0000;
        rom[5][775] = 16'h0000;
        rom[5][776] = 16'h0000;
        rom[5][777] = 16'h0000;
        rom[5][778] = 16'h0000;
        rom[5][779] = 16'h0000;
        rom[5][780] = 16'h0000;
        rom[5][781] = 16'h0000;
        rom[5][782] = 16'h0000;
        rom[5][783] = 16'h0000;
        rom[5][784] = 16'h00F5;
        rom[5][785] = 16'h0104;
        rom[5][786] = 16'h00C3;
        rom[5][787] = 16'h0082;
        rom[5][788] = 16'h01AA;
        rom[5][789] = 16'h020F;
        rom[5][790] = 16'h0186;
        rom[5][791] = 16'h015A;
        rom[5][792] = 16'h012F;
        rom[5][793] = 16'h00F5;
        rom[5][794] = 16'h00D9;
        rom[5][795] = 16'h0112;
        rom[5][796] = 16'h00BC;
        rom[5][797] = 16'h0057;
        rom[5][798] = 16'h00B4;
        rom[5][799] = 16'h013E;
        rom[5][800] = 16'h0153;
        rom[5][801] = 16'h01BF;
        rom[5][802] = 16'h0162;
        rom[5][803] = 16'h012F;
        rom[5][804] = 16'h01DC;
        rom[5][805] = 16'h01CE;
        rom[5][806] = 16'h0136;
        rom[5][807] = 16'h0104;
        rom[5][808] = 16'h01B1;
        rom[5][809] = 16'h01CE;
        rom[5][810] = 16'h0153;
        rom[5][811] = 16'h0104;
        rom[5][812] = 16'h0112;
        rom[5][813] = 16'h013E;
        rom[5][814] = 16'h0145;
        rom[5][815] = 16'h00D9;
        rom[5][816] = 16'h0000;
        rom[5][817] = 16'h0000;
        rom[5][818] = 16'h0000;
        rom[5][819] = 16'h0000;
        rom[5][820] = 16'h0000;
        rom[5][821] = 16'h0000;
        rom[5][822] = 16'h0000;
        rom[5][823] = 16'h0000;
        rom[5][824] = 16'h0000;
        rom[5][825] = 16'h0000;
        rom[5][826] = 16'h0000;
        rom[5][827] = 16'h0000;
        rom[5][828] = 16'h0000;
        rom[5][829] = 16'h0000;
        rom[5][830] = 16'h0000;
        rom[5][831] = 16'h0000;
        rom[5][832] = 16'h0000;
        rom[5][833] = 16'h0000;
        rom[5][834] = 16'h0000;
        rom[5][835] = 16'h0000;
        rom[5][836] = 16'h0000;
        rom[5][837] = 16'h0000;
        rom[5][838] = 16'h0000;
        rom[5][839] = 16'h0000;
        rom[5][840] = 16'h0000;
        rom[5][841] = 16'h0000;
        rom[5][842] = 16'h0000;
        rom[5][843] = 16'h0000;
        rom[5][844] = 16'h0000;
        rom[5][845] = 16'h0000;
        rom[5][846] = 16'h0000;
        rom[5][847] = 16'h0000;
        rom[5][848] = 16'h0000;
        rom[5][849] = 16'h0000;
        rom[5][850] = 16'h0000;
        rom[5][851] = 16'h0000;
        rom[5][852] = 16'h0000;
        rom[5][853] = 16'h0000;
        rom[5][854] = 16'h0000;
        rom[5][855] = 16'h0000;
        rom[5][856] = 16'h0000;
        rom[5][857] = 16'h0000;
        rom[5][858] = 16'h0000;
        rom[5][859] = 16'h0000;
        rom[5][860] = 16'h0000;
        rom[5][861] = 16'h0000;
        rom[5][862] = 16'h0000;
        rom[5][863] = 16'h0000;
        rom[5][864] = 16'h0000;
        rom[5][865] = 16'h0000;
        rom[5][866] = 16'h0000;
        rom[5][867] = 16'h0000;
        rom[5][868] = 16'h0000;
        rom[5][869] = 16'h0000;
        rom[5][870] = 16'h0000;
        rom[5][871] = 16'h0000;
        rom[5][872] = 16'h0000;
        rom[5][873] = 16'h0000;
        rom[5][874] = 16'h0000;
        rom[5][875] = 16'h0000;
        rom[5][876] = 16'h0000;
        rom[5][877] = 16'h0000;
        rom[5][878] = 16'h0000;
        rom[5][879] = 16'h0000;
        rom[5][880] = 16'h0000;
        rom[5][881] = 16'h0000;
        rom[5][882] = 16'hFFEA;
        rom[5][883] = 16'h007B;
        rom[5][884] = 16'h00F5;
        rom[5][885] = 16'h002B;
        rom[5][886] = 16'hFE56;
        rom[5][887] = 16'hFE4F;
        rom[5][888] = 16'hFF36;
        rom[5][889] = 16'h0090;
        rom[5][890] = 16'h0145;
        rom[5][891] = 16'h01A3;
        rom[5][892] = 16'h0194;
        rom[5][893] = 16'h0128;
        rom[5][894] = 16'h009F;
        rom[5][895] = 16'h002B;
        rom[5][896] = 16'h0033;
        rom[5][897] = 16'h002B;
        rom[5][898] = 16'hFFF2;
        rom[5][899] = 16'h0000;
        rom[5][900] = 16'h0041;
        rom[5][901] = 16'hFFF9;
        rom[5][902] = 16'h0065;
        rom[5][903] = 16'h0073;
        rom[5][904] = 16'h004F;
        rom[5][905] = 16'h0057;
        rom[5][906] = 16'h007B;
        rom[5][907] = 16'h009F;
        rom[5][908] = 16'h00A6;
        rom[5][909] = 16'h0041;
        rom[5][910] = 16'h0041;
        rom[5][911] = 16'h0057;
        rom[5][912] = 16'h0057;
        rom[5][913] = 16'h0065;
        rom[5][914] = 16'h0000;
        rom[5][915] = 16'h0000;
        rom[5][916] = 16'h0000;
        rom[5][917] = 16'h0000;
        rom[5][918] = 16'h0000;
        rom[5][919] = 16'h0000;
        rom[5][920] = 16'h0000;
        rom[5][921] = 16'h0000;
        rom[5][922] = 16'h0000;
        rom[5][923] = 16'h0000;
        rom[5][924] = 16'h0000;
        rom[5][925] = 16'h0000;
        rom[5][926] = 16'h0000;
        rom[5][927] = 16'h0000;
        rom[5][928] = 16'h0000;
        rom[5][929] = 16'h0000;
        rom[5][930] = 16'h0000;
        rom[5][931] = 16'h0000;
        rom[5][932] = 16'h0000;
        rom[5][933] = 16'h0000;
        rom[5][934] = 16'h0000;
        rom[5][935] = 16'h0000;
        rom[5][936] = 16'h0000;
        rom[5][937] = 16'h0000;
        rom[5][938] = 16'h0000;
        rom[5][939] = 16'h0000;
        rom[5][940] = 16'h0000;
        rom[5][941] = 16'h0000;
        rom[5][942] = 16'h0000;
        rom[5][943] = 16'h0000;
        rom[5][944] = 16'h0000;
        rom[5][945] = 16'h0000;
        rom[5][946] = 16'h0000;
        rom[5][947] = 16'h0000;
        rom[5][948] = 16'h0000;
        rom[5][949] = 16'h0000;
        rom[5][950] = 16'h0000;
        rom[5][951] = 16'h0000;
        rom[5][952] = 16'h0000;
        rom[5][953] = 16'h0000;
        rom[5][954] = 16'h0000;
        rom[5][955] = 16'h0000;
        rom[5][956] = 16'h0000;
        rom[5][957] = 16'h0000;
        rom[5][958] = 16'h0000;
        rom[5][959] = 16'h0000;
        rom[5][960] = 16'h0000;
        rom[5][961] = 16'h0000;
        rom[5][962] = 16'h0000;
        rom[5][963] = 16'h0000;
        rom[5][964] = 16'h0000;
        rom[5][965] = 16'h0000;
        rom[5][966] = 16'h0000;
        rom[5][967] = 16'h0000;
        rom[5][968] = 16'h0000;
        rom[5][969] = 16'h0000;
        rom[5][970] = 16'h0000;
        rom[5][971] = 16'h0000;
        rom[5][972] = 16'h0000;
        rom[5][973] = 16'h0000;
        rom[5][974] = 16'h0000;
        rom[5][975] = 16'h0000;
        rom[5][976] = 16'h0000;
        rom[5][977] = 16'h0000;
        rom[5][978] = 16'h0000;
        rom[5][979] = 16'h0000;
        rom[5][980] = 16'hFFDC;
        rom[5][981] = 16'h005E;
        rom[5][982] = 16'h00E7;
        rom[5][983] = 16'h0073;
        rom[5][984] = 16'h005E;
        rom[5][985] = 16'h00AD;
        rom[5][986] = 16'h018D;
        rom[5][987] = 16'h0119;
        rom[5][988] = 16'h0041;
        rom[5][989] = 16'h000E;
        rom[5][990] = 16'hFFE3;
        rom[5][991] = 16'hFFBF;
        rom[5][992] = 16'h009F;
        rom[5][993] = 16'h0119;
        rom[5][994] = 16'h00C3;
        rom[5][995] = 16'h00E0;
        rom[5][996] = 16'h00EE;
        rom[5][997] = 16'h00F5;
        rom[5][998] = 16'h0162;
        rom[5][999] = 16'h0170;
        rom[5][1000] = 16'h00FD;
        rom[5][1001] = 16'h0136;
        rom[5][1002] = 16'h0170;
        rom[5][1003] = 16'h013E;
        rom[5][1004] = 16'h0119;
        rom[5][1005] = 16'h00D1;
        rom[5][1006] = 16'h00E0;
        rom[5][1007] = 16'h009F;
        rom[5][1008] = 16'h00C3;
        rom[5][1009] = 16'h0065;
        rom[5][1010] = 16'h0024;
        rom[5][1011] = 16'hFFD5;
        rom[5][1012] = 16'h0000;
        rom[5][1013] = 16'h0000;
        rom[5][1014] = 16'h0000;
        rom[5][1015] = 16'h0000;
        rom[5][1016] = 16'h0000;
        rom[5][1017] = 16'h0000;
        rom[5][1018] = 16'h0000;
        rom[5][1019] = 16'h0000;
        rom[5][1020] = 16'h0000;
        rom[5][1021] = 16'h0000;
        rom[5][1022] = 16'h0000;
        rom[5][1023] = 16'h0000;
        rom[5][1024] = 16'h0000;
        rom[5][1025] = 16'h0000;
        rom[5][1026] = 16'h0000;
        rom[5][1027] = 16'h0000;
        rom[5][1028] = 16'h0000;
        rom[5][1029] = 16'h0000;
        rom[5][1030] = 16'h0000;
        rom[5][1031] = 16'h0000;
        rom[5][1032] = 16'h0000;
        rom[5][1033] = 16'h0000;
        rom[5][1034] = 16'h0000;
        rom[5][1035] = 16'h0000;
        rom[5][1036] = 16'h0000;
        rom[5][1037] = 16'h0000;
        rom[5][1038] = 16'h0000;
        rom[5][1039] = 16'h0000;
        rom[5][1040] = 16'h0000;
        rom[5][1041] = 16'h0000;
        rom[5][1042] = 16'h0000;
        rom[5][1043] = 16'h0000;
        rom[5][1044] = 16'h0000;
        rom[5][1045] = 16'h0000;
        rom[5][1046] = 16'h0000;
        rom[5][1047] = 16'h0000;
        rom[5][1048] = 16'h0000;
        rom[5][1049] = 16'h0000;
        rom[5][1050] = 16'h0000;
        rom[5][1051] = 16'h0000;
        rom[5][1052] = 16'h0000;
        rom[5][1053] = 16'h0000;
        rom[5][1054] = 16'h0000;
        rom[5][1055] = 16'h0000;
        rom[5][1056] = 16'h0000;
        rom[5][1057] = 16'h0000;
        rom[5][1058] = 16'h0000;
        rom[5][1059] = 16'h0000;
        rom[5][1060] = 16'h0000;
        rom[5][1061] = 16'h0000;
        rom[5][1062] = 16'h0000;
        rom[5][1063] = 16'h0000;
        rom[5][1064] = 16'h0000;
        rom[5][1065] = 16'h0000;
        rom[5][1066] = 16'h0000;
        rom[5][1067] = 16'h0000;
        rom[5][1068] = 16'h0000;
        rom[5][1069] = 16'h0000;
        rom[5][1070] = 16'h0000;
        rom[5][1071] = 16'h0000;
        rom[5][1072] = 16'h0000;
        rom[5][1073] = 16'h0000;
        rom[5][1074] = 16'h0000;
        rom[5][1075] = 16'h0000;
        rom[5][1076] = 16'h0000;
        rom[5][1077] = 16'h0000;
        rom[5][1078] = 16'h0041;
        rom[5][1079] = 16'h0000;
        rom[5][1080] = 16'hFFA2;
        rom[5][1081] = 16'h0000;
        rom[5][1082] = 16'h00B4;
        rom[5][1083] = 16'hFF4C;
        rom[5][1084] = 16'hFF36;
        rom[5][1085] = 16'h005E;
        rom[5][1086] = 16'h012F;
        rom[5][1087] = 16'h013E;
        rom[5][1088] = 16'h0162;
        rom[5][1089] = 16'h0136;
        rom[5][1090] = 16'h00EE;
        rom[5][1091] = 16'h0128;
        rom[5][1092] = 16'h00BC;
        rom[5][1093] = 16'h003A;
        rom[5][1094] = 16'h0073;
        rom[5][1095] = 16'h0089;
        rom[5][1096] = 16'h00B4;
        rom[5][1097] = 16'h0112;
        rom[5][1098] = 16'h00D9;
        rom[5][1099] = 16'h00CA;
        rom[5][1100] = 16'h00C3;
        rom[5][1101] = 16'h00E0;
        rom[5][1102] = 16'h00EE;
        rom[5][1103] = 16'h0082;
        rom[5][1104] = 16'h005E;
        rom[5][1105] = 16'h0016;
        rom[5][1106] = 16'hFFE3;
        rom[5][1107] = 16'hFFB8;
        rom[5][1108] = 16'hFF9B;
        rom[5][1109] = 16'hFF94;
        rom[5][1110] = 16'h0000;
        rom[5][1111] = 16'h0000;
        rom[5][1112] = 16'h0000;
        rom[5][1113] = 16'h0000;
        rom[5][1114] = 16'h0000;
        rom[5][1115] = 16'h0000;
        rom[5][1116] = 16'h0000;
        rom[5][1117] = 16'h0000;
        rom[5][1118] = 16'h0000;
        rom[5][1119] = 16'h0000;
        rom[5][1120] = 16'h0000;
        rom[5][1121] = 16'h0000;
        rom[5][1122] = 16'h0000;
        rom[5][1123] = 16'h0000;
        rom[5][1124] = 16'h0000;
        rom[5][1125] = 16'h0000;
        rom[5][1126] = 16'h0000;
        rom[5][1127] = 16'h0000;
        rom[5][1128] = 16'h0000;
        rom[5][1129] = 16'h0000;
        rom[5][1130] = 16'h0000;
        rom[5][1131] = 16'h0000;
        rom[5][1132] = 16'h0000;
        rom[5][1133] = 16'h0000;
        rom[5][1134] = 16'h0000;
        rom[5][1135] = 16'h0000;
        rom[5][1136] = 16'h0000;
        rom[5][1137] = 16'h0000;
        rom[5][1138] = 16'h0000;
        rom[5][1139] = 16'h0000;
        rom[5][1140] = 16'h0000;
        rom[5][1141] = 16'h0000;
        rom[5][1142] = 16'h0000;
        rom[5][1143] = 16'h0000;
        rom[5][1144] = 16'h0000;
        rom[5][1145] = 16'h0000;
        rom[5][1146] = 16'h0000;
        rom[5][1147] = 16'h0000;
        rom[5][1148] = 16'h0000;
        rom[5][1149] = 16'h0000;
        rom[5][1150] = 16'h0000;
        rom[5][1151] = 16'h0000;
        rom[5][1152] = 16'h0000;
        rom[5][1153] = 16'h0000;
        rom[5][1154] = 16'h0000;
        rom[5][1155] = 16'h0000;
        rom[5][1156] = 16'h0000;
        rom[5][1157] = 16'h0000;
        rom[5][1158] = 16'h0000;
        rom[5][1159] = 16'h0000;
        rom[5][1160] = 16'h0000;
        rom[5][1161] = 16'h0000;
        rom[5][1162] = 16'h0000;
        rom[5][1163] = 16'h0000;
        rom[5][1164] = 16'h0000;
        rom[5][1165] = 16'h0000;
        rom[5][1166] = 16'h0000;
        rom[5][1167] = 16'h0000;
        rom[5][1168] = 16'h0000;
        rom[5][1169] = 16'h0000;
        rom[5][1170] = 16'h0000;
        rom[5][1171] = 16'h0000;
        rom[5][1172] = 16'h0000;
        rom[5][1173] = 16'h0000;
        rom[5][1174] = 16'h0000;
        rom[5][1175] = 16'h0000;
        rom[5][1176] = 16'h00C3;
        rom[5][1177] = 16'h007B;
        rom[5][1178] = 16'h007B;
        rom[5][1179] = 16'h00BC;
        rom[5][1180] = 16'h0128;
        rom[5][1181] = 16'h01F2;
        rom[5][1182] = 16'h01BF;
        rom[5][1183] = 16'h00FD;
        rom[5][1184] = 16'h010B;
        rom[5][1185] = 16'h0169;
        rom[5][1186] = 16'h017F;
        rom[5][1187] = 16'h019B;
        rom[5][1188] = 16'h0170;
        rom[5][1189] = 16'h01CE;
        rom[5][1190] = 16'h01F2;
        rom[5][1191] = 16'h019B;
        rom[5][1192] = 16'h015A;
        rom[5][1193] = 16'h01A3;
        rom[5][1194] = 16'h01CE;
        rom[5][1195] = 16'h019B;
        rom[5][1196] = 16'h01F2;
        rom[5][1197] = 16'h013E;
        rom[5][1198] = 16'h00F5;
        rom[5][1199] = 16'h014C;
        rom[5][1200] = 16'h0145;
        rom[5][1201] = 16'h015A;
        rom[5][1202] = 16'h0121;
        rom[5][1203] = 16'h005E;
        rom[5][1204] = 16'h004F;
        rom[5][1205] = 16'h0090;
        rom[5][1206] = 16'h0098;
        rom[5][1207] = 16'h010B;
        rom[5][1208] = 16'h0000;
        rom[5][1209] = 16'h0000;
        rom[5][1210] = 16'h0000;
        rom[5][1211] = 16'h0000;
        rom[5][1212] = 16'h0000;
        rom[5][1213] = 16'h0000;
        rom[5][1214] = 16'h0000;
        rom[5][1215] = 16'h0000;
        rom[5][1216] = 16'h0000;
        rom[5][1217] = 16'h0000;
        rom[5][1218] = 16'h0000;
        rom[5][1219] = 16'h0000;
        rom[5][1220] = 16'h0000;
        rom[5][1221] = 16'h0000;
        rom[5][1222] = 16'h0000;
        rom[5][1223] = 16'h0000;
        rom[5][1224] = 16'h0000;
        rom[5][1225] = 16'h0000;
        rom[5][1226] = 16'h0000;
        rom[5][1227] = 16'h0000;
        rom[5][1228] = 16'h0000;
        rom[5][1229] = 16'h0000;
        rom[5][1230] = 16'h0000;
        rom[5][1231] = 16'h0000;
        rom[5][1232] = 16'h0000;
        rom[5][1233] = 16'h0000;
        rom[5][1234] = 16'h0000;
        rom[5][1235] = 16'h0000;
        rom[5][1236] = 16'h0000;
        rom[5][1237] = 16'h0000;
        rom[5][1238] = 16'h0000;
        rom[5][1239] = 16'h0000;
        rom[5][1240] = 16'h0000;
        rom[5][1241] = 16'h0000;
        rom[5][1242] = 16'h0000;
        rom[5][1243] = 16'h0000;
        rom[5][1244] = 16'h0000;
        rom[5][1245] = 16'h0000;
        rom[5][1246] = 16'h0000;
        rom[5][1247] = 16'h0000;
        rom[5][1248] = 16'h0000;
        rom[5][1249] = 16'h0000;
        rom[5][1250] = 16'h0000;
        rom[5][1251] = 16'h0000;
        rom[5][1252] = 16'h0000;
        rom[5][1253] = 16'h0000;
        rom[5][1254] = 16'h0000;
        rom[5][1255] = 16'h0000;
        rom[5][1256] = 16'h0000;
        rom[5][1257] = 16'h0000;
        rom[5][1258] = 16'h0000;
        rom[5][1259] = 16'h0000;
        rom[5][1260] = 16'h0000;
        rom[5][1261] = 16'h0000;
        rom[5][1262] = 16'h0000;
        rom[5][1263] = 16'h0000;
        rom[5][1264] = 16'h0000;
        rom[5][1265] = 16'h0000;
        rom[5][1266] = 16'h0000;
        rom[5][1267] = 16'h0000;
        rom[5][1268] = 16'h0000;
        rom[5][1269] = 16'h0000;
        rom[5][1270] = 16'h0000;
        rom[5][1271] = 16'h0000;
        rom[5][1272] = 16'h0000;
        rom[5][1273] = 16'h0000;
        rom[6][0] = 16'h02EF;
        rom[6][1] = 16'h02D9;
        rom[6][2] = 16'h02EF;
        rom[6][3] = 16'h02C3;
        rom[6][4] = 16'h023A;
        rom[6][5] = 16'h017F;
        rom[6][6] = 16'h00FD;
        rom[6][7] = 16'h005E;
        rom[6][8] = 16'h0065;
        rom[6][9] = 16'h010B;
        rom[6][10] = 16'h012F;
        rom[6][11] = 16'h0121;
        rom[6][12] = 16'h0119;
        rom[6][13] = 16'h0119;
        rom[6][14] = 16'h012F;
        rom[6][15] = 16'h013E;
        rom[6][16] = 16'h0112;
        rom[6][17] = 16'h00EE;
        rom[6][18] = 16'h0177;
        rom[6][19] = 16'h01AA;
        rom[6][20] = 16'h0186;
        rom[6][21] = 16'h013E;
        rom[6][22] = 16'h00EE;
        rom[6][23] = 16'h007B;
        rom[6][24] = 16'h003A;
        rom[6][25] = 16'h00CA;
        rom[6][26] = 16'h00E7;
        rom[6][27] = 16'h007B;
        rom[6][28] = 16'hFFB8;
        rom[6][29] = 16'hFFCD;
        rom[6][30] = 16'h007B;
        rom[6][31] = 16'h00C3;
        rom[6][32] = 16'h0000;
        rom[6][33] = 16'h0000;
        rom[6][34] = 16'h0000;
        rom[6][35] = 16'h0000;
        rom[6][36] = 16'h0000;
        rom[6][37] = 16'h0000;
        rom[6][38] = 16'h0000;
        rom[6][39] = 16'h0000;
        rom[6][40] = 16'h0000;
        rom[6][41] = 16'h0000;
        rom[6][42] = 16'h0000;
        rom[6][43] = 16'h0000;
        rom[6][44] = 16'h0000;
        rom[6][45] = 16'h0000;
        rom[6][46] = 16'h0000;
        rom[6][47] = 16'h0000;
        rom[6][48] = 16'h0000;
        rom[6][49] = 16'h0000;
        rom[6][50] = 16'h0000;
        rom[6][51] = 16'h0000;
        rom[6][52] = 16'h0000;
        rom[6][53] = 16'h0000;
        rom[6][54] = 16'h0000;
        rom[6][55] = 16'h0000;
        rom[6][56] = 16'h0000;
        rom[6][57] = 16'h0000;
        rom[6][58] = 16'h0000;
        rom[6][59] = 16'h0000;
        rom[6][60] = 16'h0000;
        rom[6][61] = 16'h0000;
        rom[6][62] = 16'h0000;
        rom[6][63] = 16'h0000;
        rom[6][64] = 16'h0000;
        rom[6][65] = 16'h0000;
        rom[6][66] = 16'h0000;
        rom[6][67] = 16'h0000;
        rom[6][68] = 16'h0000;
        rom[6][69] = 16'h0000;
        rom[6][70] = 16'h0000;
        rom[6][71] = 16'h0000;
        rom[6][72] = 16'h0000;
        rom[6][73] = 16'h0000;
        rom[6][74] = 16'h0000;
        rom[6][75] = 16'h0000;
        rom[6][76] = 16'h0000;
        rom[6][77] = 16'h0000;
        rom[6][78] = 16'h0000;
        rom[6][79] = 16'h0000;
        rom[6][80] = 16'h0000;
        rom[6][81] = 16'h0000;
        rom[6][82] = 16'h0000;
        rom[6][83] = 16'h0000;
        rom[6][84] = 16'h0000;
        rom[6][85] = 16'h0000;
        rom[6][86] = 16'h0000;
        rom[6][87] = 16'h0000;
        rom[6][88] = 16'h0000;
        rom[6][89] = 16'h0000;
        rom[6][90] = 16'h0000;
        rom[6][91] = 16'h0000;
        rom[6][92] = 16'h0000;
        rom[6][93] = 16'h0000;
        rom[6][94] = 16'h0000;
        rom[6][95] = 16'h0000;
        rom[6][96] = 16'h0000;
        rom[6][97] = 16'h0000;
        rom[6][98] = 16'h00F5;
        rom[6][99] = 16'h00EE;
        rom[6][100] = 16'h0119;
        rom[6][101] = 16'h00C3;
        rom[6][102] = 16'h00D1;
        rom[6][103] = 16'h0186;
        rom[6][104] = 16'h019B;
        rom[6][105] = 16'h0128;
        rom[6][106] = 16'h0033;
        rom[6][107] = 16'h004F;
        rom[6][108] = 16'h0073;
        rom[6][109] = 16'h007B;
        rom[6][110] = 16'h0073;
        rom[6][111] = 16'h0057;
        rom[6][112] = 16'h0057;
        rom[6][113] = 16'h007B;
        rom[6][114] = 16'h00B4;
        rom[6][115] = 16'h00C3;
        rom[6][116] = 16'hFFEA;
        rom[6][117] = 16'hFF7E;
        rom[6][118] = 16'hFF44;
        rom[6][119] = 16'hFEFC;
        rom[6][120] = 16'hFEFC;
        rom[6][121] = 16'hFF4C;
        rom[6][122] = 16'hFF5A;
        rom[6][123] = 16'hFFA9;
        rom[6][124] = 16'hFFC6;
        rom[6][125] = 16'hFFBF;
        rom[6][126] = 16'hFF70;
        rom[6][127] = 16'hFF03;
        rom[6][128] = 16'hFE9E;
        rom[6][129] = 16'hFE39;
        rom[6][130] = 16'h0000;
        rom[6][131] = 16'h0000;
        rom[6][132] = 16'h0000;
        rom[6][133] = 16'h0000;
        rom[6][134] = 16'h0000;
        rom[6][135] = 16'h0000;
        rom[6][136] = 16'h0000;
        rom[6][137] = 16'h0000;
        rom[6][138] = 16'h0000;
        rom[6][139] = 16'h0000;
        rom[6][140] = 16'h0000;
        rom[6][141] = 16'h0000;
        rom[6][142] = 16'h0000;
        rom[6][143] = 16'h0000;
        rom[6][144] = 16'h0000;
        rom[6][145] = 16'h0000;
        rom[6][146] = 16'h0000;
        rom[6][147] = 16'h0000;
        rom[6][148] = 16'h0000;
        rom[6][149] = 16'h0000;
        rom[6][150] = 16'h0000;
        rom[6][151] = 16'h0000;
        rom[6][152] = 16'h0000;
        rom[6][153] = 16'h0000;
        rom[6][154] = 16'h0000;
        rom[6][155] = 16'h0000;
        rom[6][156] = 16'h0000;
        rom[6][157] = 16'h0000;
        rom[6][158] = 16'h0000;
        rom[6][159] = 16'h0000;
        rom[6][160] = 16'h0000;
        rom[6][161] = 16'h0000;
        rom[6][162] = 16'h0000;
        rom[6][163] = 16'h0000;
        rom[6][164] = 16'h0000;
        rom[6][165] = 16'h0000;
        rom[6][166] = 16'h0000;
        rom[6][167] = 16'h0000;
        rom[6][168] = 16'h0000;
        rom[6][169] = 16'h0000;
        rom[6][170] = 16'h0000;
        rom[6][171] = 16'h0000;
        rom[6][172] = 16'h0000;
        rom[6][173] = 16'h0000;
        rom[6][174] = 16'h0000;
        rom[6][175] = 16'h0000;
        rom[6][176] = 16'h0000;
        rom[6][177] = 16'h0000;
        rom[6][178] = 16'h0000;
        rom[6][179] = 16'h0000;
        rom[6][180] = 16'h0000;
        rom[6][181] = 16'h0000;
        rom[6][182] = 16'h0000;
        rom[6][183] = 16'h0000;
        rom[6][184] = 16'h0000;
        rom[6][185] = 16'h0000;
        rom[6][186] = 16'h0000;
        rom[6][187] = 16'h0000;
        rom[6][188] = 16'h0000;
        rom[6][189] = 16'h0000;
        rom[6][190] = 16'h0000;
        rom[6][191] = 16'h0000;
        rom[6][192] = 16'h0000;
        rom[6][193] = 16'h0000;
        rom[6][194] = 16'h0000;
        rom[6][195] = 16'h0000;
        rom[6][196] = 16'h0089;
        rom[6][197] = 16'hFFCD;
        rom[6][198] = 16'hFF61;
        rom[6][199] = 16'hFEEE;
        rom[6][200] = 16'hFED1;
        rom[6][201] = 16'hFEB4;
        rom[6][202] = 16'hFF27;
        rom[6][203] = 16'h004F;
        rom[6][204] = 16'hFFB1;
        rom[6][205] = 16'hFEA6;
        rom[6][206] = 16'hFE56;
        rom[6][207] = 16'hFE4F;
        rom[6][208] = 16'hFE56;
        rom[6][209] = 16'hFE48;
        rom[6][210] = 16'hFE7A;
        rom[6][211] = 16'hFEAD;
        rom[6][212] = 16'hFE97;
        rom[6][213] = 16'hFEE7;
        rom[6][214] = 16'hFF12;
        rom[6][215] = 16'hFF12;
        rom[6][216] = 16'hFF0B;
        rom[6][217] = 16'hFE97;
        rom[6][218] = 16'hFDE3;
        rom[6][219] = 16'hFD2E;
        rom[6][220] = 16'hFD0A;
        rom[6][221] = 16'h0378;
        rom[6][222] = 16'h035B;
        rom[6][223] = 16'hFCD8;
        rom[6][224] = 16'hFEAD;
        rom[6][225] = 16'hFEAD;
        rom[6][226] = 16'hFCC2;
        rom[6][227] = 16'h031A;
        rom[6][228] = 16'h0000;
        rom[6][229] = 16'h0000;
        rom[6][230] = 16'h0000;
        rom[6][231] = 16'h0000;
        rom[6][232] = 16'h0000;
        rom[6][233] = 16'h0000;
        rom[6][234] = 16'h0000;
        rom[6][235] = 16'h0000;
        rom[6][236] = 16'h0000;
        rom[6][237] = 16'h0000;
        rom[6][238] = 16'h0000;
        rom[6][239] = 16'h0000;
        rom[6][240] = 16'h0000;
        rom[6][241] = 16'h0000;
        rom[6][242] = 16'h0000;
        rom[6][243] = 16'h0000;
        rom[6][244] = 16'h0000;
        rom[6][245] = 16'h0000;
        rom[6][246] = 16'h0000;
        rom[6][247] = 16'h0000;
        rom[6][248] = 16'h0000;
        rom[6][249] = 16'h0000;
        rom[6][250] = 16'h0000;
        rom[6][251] = 16'h0000;
        rom[6][252] = 16'h0000;
        rom[6][253] = 16'h0000;
        rom[6][254] = 16'h0000;
        rom[6][255] = 16'h0000;
        rom[6][256] = 16'h0000;
        rom[6][257] = 16'h0000;
        rom[6][258] = 16'h0000;
        rom[6][259] = 16'h0000;
        rom[6][260] = 16'h0000;
        rom[6][261] = 16'h0000;
        rom[6][262] = 16'h0000;
        rom[6][263] = 16'h0000;
        rom[6][264] = 16'h0000;
        rom[6][265] = 16'h0000;
        rom[6][266] = 16'h0000;
        rom[6][267] = 16'h0000;
        rom[6][268] = 16'h0000;
        rom[6][269] = 16'h0000;
        rom[6][270] = 16'h0000;
        rom[6][271] = 16'h0000;
        rom[6][272] = 16'h0000;
        rom[6][273] = 16'h0000;
        rom[6][274] = 16'h0000;
        rom[6][275] = 16'h0000;
        rom[6][276] = 16'h0000;
        rom[6][277] = 16'h0000;
        rom[6][278] = 16'h0000;
        rom[6][279] = 16'h0000;
        rom[6][280] = 16'h0000;
        rom[6][281] = 16'h0000;
        rom[6][282] = 16'h0000;
        rom[6][283] = 16'h0000;
        rom[6][284] = 16'h0000;
        rom[6][285] = 16'h0000;
        rom[6][286] = 16'h0000;
        rom[6][287] = 16'h0000;
        rom[6][288] = 16'h0000;
        rom[6][289] = 16'h0000;
        rom[6][290] = 16'h0000;
        rom[6][291] = 16'h0000;
        rom[6][292] = 16'h0000;
        rom[6][293] = 16'h0000;
        rom[6][294] = 16'h0089;
        rom[6][295] = 16'hFFE3;
        rom[6][296] = 16'hFFBF;
        rom[6][297] = 16'h005E;
        rom[6][298] = 16'h00A6;
        rom[6][299] = 16'h015A;
        rom[6][300] = 16'h0153;
        rom[6][301] = 16'h00AD;
        rom[6][302] = 16'h0104;
        rom[6][303] = 16'h014C;
        rom[6][304] = 16'h0194;
        rom[6][305] = 16'h01A3;
        rom[6][306] = 16'h01AA;
        rom[6][307] = 16'h0169;
        rom[6][308] = 16'h00E0;
        rom[6][309] = 16'h00B4;
        rom[6][310] = 16'h00BC;
        rom[6][311] = 16'h0048;
        rom[6][312] = 16'h00C3;
        rom[6][313] = 16'h00D9;
        rom[6][314] = 16'h00AD;
        rom[6][315] = 16'h0098;
        rom[6][316] = 16'h007B;
        rom[6][317] = 16'h0090;
        rom[6][318] = 16'h0065;
        rom[6][319] = 16'h009F;
        rom[6][320] = 16'h00A6;
        rom[6][321] = 16'h0073;
        rom[6][322] = 16'h0041;
        rom[6][323] = 16'h01DC;
        rom[6][324] = 16'h02D2;
        rom[6][325] = 16'h0321;
        rom[6][326] = 16'h0000;
        rom[6][327] = 16'h0000;
        rom[6][328] = 16'h0000;
        rom[6][329] = 16'h0000;
        rom[6][330] = 16'h0000;
        rom[6][331] = 16'h0000;
        rom[6][332] = 16'h0000;
        rom[6][333] = 16'h0000;
        rom[6][334] = 16'h0000;
        rom[6][335] = 16'h0000;
        rom[6][336] = 16'h0000;
        rom[6][337] = 16'h0000;
        rom[6][338] = 16'h0000;
        rom[6][339] = 16'h0000;
        rom[6][340] = 16'h0000;
        rom[6][341] = 16'h0000;
        rom[6][342] = 16'h0000;
        rom[6][343] = 16'h0000;
        rom[6][344] = 16'h0000;
        rom[6][345] = 16'h0000;
        rom[6][346] = 16'h0000;
        rom[6][347] = 16'h0000;
        rom[6][348] = 16'h0000;
        rom[6][349] = 16'h0000;
        rom[6][350] = 16'h0000;
        rom[6][351] = 16'h0000;
        rom[6][352] = 16'h0000;
        rom[6][353] = 16'h0000;
        rom[6][354] = 16'h0000;
        rom[6][355] = 16'h0000;
        rom[6][356] = 16'h0000;
        rom[6][357] = 16'h0000;
        rom[6][358] = 16'h0000;
        rom[6][359] = 16'h0000;
        rom[6][360] = 16'h0000;
        rom[6][361] = 16'h0000;
        rom[6][362] = 16'h0000;
        rom[6][363] = 16'h0000;
        rom[6][364] = 16'h0000;
        rom[6][365] = 16'h0000;
        rom[6][366] = 16'h0000;
        rom[6][367] = 16'h0000;
        rom[6][368] = 16'h0000;
        rom[6][369] = 16'h0000;
        rom[6][370] = 16'h0000;
        rom[6][371] = 16'h0000;
        rom[6][372] = 16'h0000;
        rom[6][373] = 16'h0000;
        rom[6][374] = 16'h0000;
        rom[6][375] = 16'h0000;
        rom[6][376] = 16'h0000;
        rom[6][377] = 16'h0000;
        rom[6][378] = 16'h0000;
        rom[6][379] = 16'h0000;
        rom[6][380] = 16'h0000;
        rom[6][381] = 16'h0000;
        rom[6][382] = 16'h0000;
        rom[6][383] = 16'h0000;
        rom[6][384] = 16'h0000;
        rom[6][385] = 16'h0000;
        rom[6][386] = 16'h0000;
        rom[6][387] = 16'h0000;
        rom[6][388] = 16'h0000;
        rom[6][389] = 16'h0000;
        rom[6][390] = 16'h0000;
        rom[6][391] = 16'h0000;
        rom[6][392] = 16'h015A;
        rom[6][393] = 16'h00EE;
        rom[6][394] = 16'h00BC;
        rom[6][395] = 16'h00C3;
        rom[6][396] = 16'h0090;
        rom[6][397] = 16'h0024;
        rom[6][398] = 16'h0041;
        rom[6][399] = 16'h00AD;
        rom[6][400] = 16'h00AD;
        rom[6][401] = 16'hFFCD;
        rom[6][402] = 16'hFF9B;
        rom[6][403] = 16'hFF77;
        rom[6][404] = 16'hFF70;
        rom[6][405] = 16'hFFCD;
        rom[6][406] = 16'h002B;
        rom[6][407] = 16'h0065;
        rom[6][408] = 16'h007B;
        rom[6][409] = 16'h0089;
        rom[6][410] = 16'h003A;
        rom[6][411] = 16'h001D;
        rom[6][412] = 16'h001D;
        rom[6][413] = 16'h005E;
        rom[6][414] = 16'hFFEA;
        rom[6][415] = 16'hFF68;
        rom[6][416] = 16'hFFCD;
        rom[6][417] = 16'hFF68;
        rom[6][418] = 16'hFF3D;
        rom[6][419] = 16'hFFA2;
        rom[6][420] = 16'h00D1;
        rom[6][421] = 16'hFFEA;
        rom[6][422] = 16'hFEC2;
        rom[6][423] = 16'hFEAD;
        rom[6][424] = 16'h0000;
        rom[6][425] = 16'h0000;
        rom[6][426] = 16'h0000;
        rom[6][427] = 16'h0000;
        rom[6][428] = 16'h0000;
        rom[6][429] = 16'h0000;
        rom[6][430] = 16'h0000;
        rom[6][431] = 16'h0000;
        rom[6][432] = 16'h0000;
        rom[6][433] = 16'h0000;
        rom[6][434] = 16'h0000;
        rom[6][435] = 16'h0000;
        rom[6][436] = 16'h0000;
        rom[6][437] = 16'h0000;
        rom[6][438] = 16'h0000;
        rom[6][439] = 16'h0000;
        rom[6][440] = 16'h0000;
        rom[6][441] = 16'h0000;
        rom[6][442] = 16'h0000;
        rom[6][443] = 16'h0000;
        rom[6][444] = 16'h0000;
        rom[6][445] = 16'h0000;
        rom[6][446] = 16'h0000;
        rom[6][447] = 16'h0000;
        rom[6][448] = 16'h0000;
        rom[6][449] = 16'h0000;
        rom[6][450] = 16'h0000;
        rom[6][451] = 16'h0000;
        rom[6][452] = 16'h0000;
        rom[6][453] = 16'h0000;
        rom[6][454] = 16'h0000;
        rom[6][455] = 16'h0000;
        rom[6][456] = 16'h0000;
        rom[6][457] = 16'h0000;
        rom[6][458] = 16'h0000;
        rom[6][459] = 16'h0000;
        rom[6][460] = 16'h0000;
        rom[6][461] = 16'h0000;
        rom[6][462] = 16'h0000;
        rom[6][463] = 16'h0000;
        rom[6][464] = 16'h0000;
        rom[6][465] = 16'h0000;
        rom[6][466] = 16'h0000;
        rom[6][467] = 16'h0000;
        rom[6][468] = 16'h0000;
        rom[6][469] = 16'h0000;
        rom[6][470] = 16'h0000;
        rom[6][471] = 16'h0000;
        rom[6][472] = 16'h0000;
        rom[6][473] = 16'h0000;
        rom[6][474] = 16'h0000;
        rom[6][475] = 16'h0000;
        rom[6][476] = 16'h0000;
        rom[6][477] = 16'h0000;
        rom[6][478] = 16'h0000;
        rom[6][479] = 16'h0000;
        rom[6][480] = 16'h0000;
        rom[6][481] = 16'h0000;
        rom[6][482] = 16'h0000;
        rom[6][483] = 16'h0000;
        rom[6][484] = 16'h0000;
        rom[6][485] = 16'h0000;
        rom[6][486] = 16'h0000;
        rom[6][487] = 16'h0000;
        rom[6][488] = 16'h0000;
        rom[6][489] = 16'h0000;
        rom[6][490] = 16'hFE15;
        rom[6][491] = 16'hFDCD;
        rom[6][492] = 16'hFE07;
        rom[6][493] = 16'hFE15;
        rom[6][494] = 16'hFE81;
        rom[6][495] = 16'hFEFC;
        rom[6][496] = 16'hFF7E;
        rom[6][497] = 16'h0016;
        rom[6][498] = 16'hFEFC;
        rom[6][499] = 16'hFE41;
        rom[6][500] = 16'hFE24;
        rom[6][501] = 16'hFE48;
        rom[6][502] = 16'hFE39;
        rom[6][503] = 16'hFE56;
        rom[6][504] = 16'hFE7A;
        rom[6][505] = 16'hFEAD;
        rom[6][506] = 16'hFEFC;
        rom[6][507] = 16'hFF20;
        rom[6][508] = 16'hFF12;
        rom[6][509] = 16'hFF3D;
        rom[6][510] = 16'hFF68;
        rom[6][511] = 16'hFF9B;
        rom[6][512] = 16'hFF19;
        rom[6][513] = 16'hFF12;
        rom[6][514] = 16'hFEAD;
        rom[6][515] = 16'hFE41;
        rom[6][516] = 16'hFE15;
        rom[6][517] = 16'hFDC6;
        rom[6][518] = 16'hFE15;
        rom[6][519] = 16'hFDE3;
        rom[6][520] = 16'hFED1;
        rom[6][521] = 16'hFF0B;
        rom[6][522] = 16'h0000;
        rom[6][523] = 16'h0000;
        rom[6][524] = 16'h0000;
        rom[6][525] = 16'h0000;
        rom[6][526] = 16'h0000;
        rom[6][527] = 16'h0000;
        rom[6][528] = 16'h0000;
        rom[6][529] = 16'h0000;
        rom[6][530] = 16'h0000;
        rom[6][531] = 16'h0000;
        rom[6][532] = 16'h0000;
        rom[6][533] = 16'h0000;
        rom[6][534] = 16'h0000;
        rom[6][535] = 16'h0000;
        rom[6][536] = 16'h0000;
        rom[6][537] = 16'h0000;
        rom[6][538] = 16'h0000;
        rom[6][539] = 16'h0000;
        rom[6][540] = 16'h0000;
        rom[6][541] = 16'h0000;
        rom[6][542] = 16'h0000;
        rom[6][543] = 16'h0000;
        rom[6][544] = 16'h0000;
        rom[6][545] = 16'h0000;
        rom[6][546] = 16'h0000;
        rom[6][547] = 16'h0000;
        rom[6][548] = 16'h0000;
        rom[6][549] = 16'h0000;
        rom[6][550] = 16'h0000;
        rom[6][551] = 16'h0000;
        rom[6][552] = 16'h0000;
        rom[6][553] = 16'h0000;
        rom[6][554] = 16'h0000;
        rom[6][555] = 16'h0000;
        rom[6][556] = 16'h0000;
        rom[6][557] = 16'h0000;
        rom[6][558] = 16'h0000;
        rom[6][559] = 16'h0000;
        rom[6][560] = 16'h0000;
        rom[6][561] = 16'h0000;
        rom[6][562] = 16'h0000;
        rom[6][563] = 16'h0000;
        rom[6][564] = 16'h0000;
        rom[6][565] = 16'h0000;
        rom[6][566] = 16'h0000;
        rom[6][567] = 16'h0000;
        rom[6][568] = 16'h0000;
        rom[6][569] = 16'h0000;
        rom[6][570] = 16'h0000;
        rom[6][571] = 16'h0000;
        rom[6][572] = 16'h0000;
        rom[6][573] = 16'h0000;
        rom[6][574] = 16'h0000;
        rom[6][575] = 16'h0000;
        rom[6][576] = 16'h0000;
        rom[6][577] = 16'h0000;
        rom[6][578] = 16'h0000;
        rom[6][579] = 16'h0000;
        rom[6][580] = 16'h0000;
        rom[6][581] = 16'h0000;
        rom[6][582] = 16'h0000;
        rom[6][583] = 16'h0000;
        rom[6][584] = 16'h0000;
        rom[6][585] = 16'h0000;
        rom[6][586] = 16'h0000;
        rom[6][587] = 16'h0000;
        rom[6][588] = 16'h010B;
        rom[6][589] = 16'h00E0;
        rom[6][590] = 16'h0048;
        rom[6][591] = 16'h0089;
        rom[6][592] = 16'h00E7;
        rom[6][593] = 16'h00EE;
        rom[6][594] = 16'h00E7;
        rom[6][595] = 16'h00BC;
        rom[6][596] = 16'hFF8D;
        rom[6][597] = 16'hFF5A;
        rom[6][598] = 16'hFFD5;
        rom[6][599] = 16'hFFCD;
        rom[6][600] = 16'hFF5A;
        rom[6][601] = 16'hFF12;
        rom[6][602] = 16'hFEEE;
        rom[6][603] = 16'hFF03;
        rom[6][604] = 16'hFF2F;
        rom[6][605] = 16'hFEE7;
        rom[6][606] = 16'hFF19;
        rom[6][607] = 16'hFF68;
        rom[6][608] = 16'hFF85;
        rom[6][609] = 16'hFF7E;
        rom[6][610] = 16'hFEDF;
        rom[6][611] = 16'hFE89;
        rom[6][612] = 16'hFF77;
        rom[6][613] = 16'hFF85;
        rom[6][614] = 16'hFF2F;
        rom[6][615] = 16'hFF44;
        rom[6][616] = 16'hFF0B;
        rom[6][617] = 16'h00BC;
        rom[6][618] = 16'h0024;
        rom[6][619] = 16'hFF20;
        rom[6][620] = 16'h0000;
        rom[6][621] = 16'h0000;
        rom[6][622] = 16'h0000;
        rom[6][623] = 16'h0000;
        rom[6][624] = 16'h0000;
        rom[6][625] = 16'h0000;
        rom[6][626] = 16'h0000;
        rom[6][627] = 16'h0000;
        rom[6][628] = 16'h0000;
        rom[6][629] = 16'h0000;
        rom[6][630] = 16'h0000;
        rom[6][631] = 16'h0000;
        rom[6][632] = 16'h0000;
        rom[6][633] = 16'h0000;
        rom[6][634] = 16'h0000;
        rom[6][635] = 16'h0000;
        rom[6][636] = 16'h0000;
        rom[6][637] = 16'h0000;
        rom[6][638] = 16'h0000;
        rom[6][639] = 16'h0000;
        rom[6][640] = 16'h0000;
        rom[6][641] = 16'h0000;
        rom[6][642] = 16'h0000;
        rom[6][643] = 16'h0000;
        rom[6][644] = 16'h0000;
        rom[6][645] = 16'h0000;
        rom[6][646] = 16'h0000;
        rom[6][647] = 16'h0000;
        rom[6][648] = 16'h0000;
        rom[6][649] = 16'h0000;
        rom[6][650] = 16'h0000;
        rom[6][651] = 16'h0000;
        rom[6][652] = 16'h0000;
        rom[6][653] = 16'h0000;
        rom[6][654] = 16'h0000;
        rom[6][655] = 16'h0000;
        rom[6][656] = 16'h0000;
        rom[6][657] = 16'h0000;
        rom[6][658] = 16'h0000;
        rom[6][659] = 16'h0000;
        rom[6][660] = 16'h0000;
        rom[6][661] = 16'h0000;
        rom[6][662] = 16'h0000;
        rom[6][663] = 16'h0000;
        rom[6][664] = 16'h0000;
        rom[6][665] = 16'h0000;
        rom[6][666] = 16'h0000;
        rom[6][667] = 16'h0000;
        rom[6][668] = 16'h0000;
        rom[6][669] = 16'h0000;
        rom[6][670] = 16'h0000;
        rom[6][671] = 16'h0000;
        rom[6][672] = 16'h0000;
        rom[6][673] = 16'h0000;
        rom[6][674] = 16'h0000;
        rom[6][675] = 16'h0000;
        rom[6][676] = 16'h0000;
        rom[6][677] = 16'h0000;
        rom[6][678] = 16'h0000;
        rom[6][679] = 16'h0000;
        rom[6][680] = 16'h0000;
        rom[6][681] = 16'h0000;
        rom[6][682] = 16'h0000;
        rom[6][683] = 16'h0000;
        rom[6][684] = 16'h0000;
        rom[6][685] = 16'h0000;
        rom[6][686] = 16'hFCE6;
        rom[6][687] = 16'hFD2E;
        rom[6][688] = 16'hFD52;
        rom[6][689] = 16'hFDB7;
        rom[6][690] = 16'hFE00;
        rom[6][691] = 16'hFE65;
        rom[6][692] = 16'hFEA6;
        rom[6][693] = 16'hFF53;
        rom[6][694] = 16'hFEBB;
        rom[6][695] = 16'hFD9B;
        rom[6][696] = 16'hFD61;
        rom[6][697] = 16'hFDDB;
        rom[6][698] = 16'hFE39;
        rom[6][699] = 16'hFE4F;
        rom[6][700] = 16'hFE41;
        rom[6][701] = 16'hFDD4;
        rom[6][702] = 16'hFDA9;
        rom[6][703] = 16'hFE41;
        rom[6][704] = 16'hFFD5;
        rom[6][705] = 16'h007B;
        rom[6][706] = 16'h006C;
        rom[6][707] = 16'h0048;
        rom[6][708] = 16'hFFDC;
        rom[6][709] = 16'hFF8D;
        rom[6][710] = 16'hFFDC;
        rom[6][711] = 16'hFF44;
        rom[6][712] = 16'hFF53;
        rom[6][713] = 16'hFFA2;
        rom[6][714] = 16'h001D;
        rom[6][715] = 16'hFFDC;
        rom[6][716] = 16'hFFC6;
        rom[6][717] = 16'h0007;
        rom[6][718] = 16'h0000;
        rom[6][719] = 16'h0000;
        rom[6][720] = 16'h0000;
        rom[6][721] = 16'h0000;
        rom[6][722] = 16'h0000;
        rom[6][723] = 16'h0000;
        rom[6][724] = 16'h0000;
        rom[6][725] = 16'h0000;
        rom[6][726] = 16'h0000;
        rom[6][727] = 16'h0000;
        rom[6][728] = 16'h0000;
        rom[6][729] = 16'h0000;
        rom[6][730] = 16'h0000;
        rom[6][731] = 16'h0000;
        rom[6][732] = 16'h0000;
        rom[6][733] = 16'h0000;
        rom[6][734] = 16'h0000;
        rom[6][735] = 16'h0000;
        rom[6][736] = 16'h0000;
        rom[6][737] = 16'h0000;
        rom[6][738] = 16'h0000;
        rom[6][739] = 16'h0000;
        rom[6][740] = 16'h0000;
        rom[6][741] = 16'h0000;
        rom[6][742] = 16'h0000;
        rom[6][743] = 16'h0000;
        rom[6][744] = 16'h0000;
        rom[6][745] = 16'h0000;
        rom[6][746] = 16'h0000;
        rom[6][747] = 16'h0000;
        rom[6][748] = 16'h0000;
        rom[6][749] = 16'h0000;
        rom[6][750] = 16'h0000;
        rom[6][751] = 16'h0000;
        rom[6][752] = 16'h0000;
        rom[6][753] = 16'h0000;
        rom[6][754] = 16'h0000;
        rom[6][755] = 16'h0000;
        rom[6][756] = 16'h0000;
        rom[6][757] = 16'h0000;
        rom[6][758] = 16'h0000;
        rom[6][759] = 16'h0000;
        rom[6][760] = 16'h0000;
        rom[6][761] = 16'h0000;
        rom[6][762] = 16'h0000;
        rom[6][763] = 16'h0000;
        rom[6][764] = 16'h0000;
        rom[6][765] = 16'h0000;
        rom[6][766] = 16'h0000;
        rom[6][767] = 16'h0000;
        rom[6][768] = 16'h0000;
        rom[6][769] = 16'h0000;
        rom[6][770] = 16'h0000;
        rom[6][771] = 16'h0000;
        rom[6][772] = 16'h0000;
        rom[6][773] = 16'h0000;
        rom[6][774] = 16'h0000;
        rom[6][775] = 16'h0000;
        rom[6][776] = 16'h0000;
        rom[6][777] = 16'h0000;
        rom[6][778] = 16'h0000;
        rom[6][779] = 16'h0000;
        rom[6][780] = 16'h0000;
        rom[6][781] = 16'h0000;
        rom[6][782] = 16'h0000;
        rom[6][783] = 16'h0000;
        rom[6][784] = 16'hFEF5;
        rom[6][785] = 16'hFF20;
        rom[6][786] = 16'hFFB8;
        rom[6][787] = 16'h004F;
        rom[6][788] = 16'hFFEA;
        rom[6][789] = 16'hFF77;
        rom[6][790] = 16'hFF5A;
        rom[6][791] = 16'hFF20;
        rom[6][792] = 16'hFF8D;
        rom[6][793] = 16'hFFEA;
        rom[6][794] = 16'h00E7;
        rom[6][795] = 16'h0170;
        rom[6][796] = 16'h0153;
        rom[6][797] = 16'h0177;
        rom[6][798] = 16'h01BF;
        rom[6][799] = 16'h01F9;
        rom[6][800] = 16'h0241;
        rom[6][801] = 16'h02C3;
        rom[6][802] = 16'h020F;
        rom[6][803] = 16'h0186;
        rom[6][804] = 16'h00FD;
        rom[6][805] = 16'h00BC;
        rom[6][806] = 16'h00A6;
        rom[6][807] = 16'h0112;
        rom[6][808] = 16'h0104;
        rom[6][809] = 16'h0082;
        rom[6][810] = 16'hFFE3;
        rom[6][811] = 16'hFF8D;
        rom[6][812] = 16'hFFA9;
        rom[6][813] = 16'hFFEA;
        rom[6][814] = 16'h00CA;
        rom[6][815] = 16'h0089;
        rom[6][816] = 16'h0000;
        rom[6][817] = 16'h0000;
        rom[6][818] = 16'h0000;
        rom[6][819] = 16'h0000;
        rom[6][820] = 16'h0000;
        rom[6][821] = 16'h0000;
        rom[6][822] = 16'h0000;
        rom[6][823] = 16'h0000;
        rom[6][824] = 16'h0000;
        rom[6][825] = 16'h0000;
        rom[6][826] = 16'h0000;
        rom[6][827] = 16'h0000;
        rom[6][828] = 16'h0000;
        rom[6][829] = 16'h0000;
        rom[6][830] = 16'h0000;
        rom[6][831] = 16'h0000;
        rom[6][832] = 16'h0000;
        rom[6][833] = 16'h0000;
        rom[6][834] = 16'h0000;
        rom[6][835] = 16'h0000;
        rom[6][836] = 16'h0000;
        rom[6][837] = 16'h0000;
        rom[6][838] = 16'h0000;
        rom[6][839] = 16'h0000;
        rom[6][840] = 16'h0000;
        rom[6][841] = 16'h0000;
        rom[6][842] = 16'h0000;
        rom[6][843] = 16'h0000;
        rom[6][844] = 16'h0000;
        rom[6][845] = 16'h0000;
        rom[6][846] = 16'h0000;
        rom[6][847] = 16'h0000;
        rom[6][848] = 16'h0000;
        rom[6][849] = 16'h0000;
        rom[6][850] = 16'h0000;
        rom[6][851] = 16'h0000;
        rom[6][852] = 16'h0000;
        rom[6][853] = 16'h0000;
        rom[6][854] = 16'h0000;
        rom[6][855] = 16'h0000;
        rom[6][856] = 16'h0000;
        rom[6][857] = 16'h0000;
        rom[6][858] = 16'h0000;
        rom[6][859] = 16'h0000;
        rom[6][860] = 16'h0000;
        rom[6][861] = 16'h0000;
        rom[6][862] = 16'h0000;
        rom[6][863] = 16'h0000;
        rom[6][864] = 16'h0000;
        rom[6][865] = 16'h0000;
        rom[6][866] = 16'h0000;
        rom[6][867] = 16'h0000;
        rom[6][868] = 16'h0000;
        rom[6][869] = 16'h0000;
        rom[6][870] = 16'h0000;
        rom[6][871] = 16'h0000;
        rom[6][872] = 16'h0000;
        rom[6][873] = 16'h0000;
        rom[6][874] = 16'h0000;
        rom[6][875] = 16'h0000;
        rom[6][876] = 16'h0000;
        rom[6][877] = 16'h0000;
        rom[6][878] = 16'h0000;
        rom[6][879] = 16'h0000;
        rom[6][880] = 16'h0000;
        rom[6][881] = 16'h0000;
        rom[6][882] = 16'h004F;
        rom[6][883] = 16'h0121;
        rom[6][884] = 16'h00A6;
        rom[6][885] = 16'h0016;
        rom[6][886] = 16'hFEE7;
        rom[6][887] = 16'hFDD4;
        rom[6][888] = 16'hFEC2;
        rom[6][889] = 16'hFF12;
        rom[6][890] = 16'h00A6;
        rom[6][891] = 16'h005E;
        rom[6][892] = 16'hFFF9;
        rom[6][893] = 16'hFFB1;
        rom[6][894] = 16'hFF61;
        rom[6][895] = 16'hFF36;
        rom[6][896] = 16'hFF36;
        rom[6][897] = 16'hFEE7;
        rom[6][898] = 16'hFEDF;
        rom[6][899] = 16'hFE41;
        rom[6][900] = 16'hFEA6;
        rom[6][901] = 16'hFF0B;
        rom[6][902] = 16'hFF4C;
        rom[6][903] = 16'hFF7E;
        rom[6][904] = 16'hFF68;
        rom[6][905] = 16'hFF5A;
        rom[6][906] = 16'hFF7E;
        rom[6][907] = 16'hFF0B;
        rom[6][908] = 16'hFE9E;
        rom[6][909] = 16'hFE5D;
        rom[6][910] = 16'hFE7A;
        rom[6][911] = 16'hFE90;
        rom[6][912] = 16'hFE56;
        rom[6][913] = 16'hFEAD;
        rom[6][914] = 16'h0000;
        rom[6][915] = 16'h0000;
        rom[6][916] = 16'h0000;
        rom[6][917] = 16'h0000;
        rom[6][918] = 16'h0000;
        rom[6][919] = 16'h0000;
        rom[6][920] = 16'h0000;
        rom[6][921] = 16'h0000;
        rom[6][922] = 16'h0000;
        rom[6][923] = 16'h0000;
        rom[6][924] = 16'h0000;
        rom[6][925] = 16'h0000;
        rom[6][926] = 16'h0000;
        rom[6][927] = 16'h0000;
        rom[6][928] = 16'h0000;
        rom[6][929] = 16'h0000;
        rom[6][930] = 16'h0000;
        rom[6][931] = 16'h0000;
        rom[6][932] = 16'h0000;
        rom[6][933] = 16'h0000;
        rom[6][934] = 16'h0000;
        rom[6][935] = 16'h0000;
        rom[6][936] = 16'h0000;
        rom[6][937] = 16'h0000;
        rom[6][938] = 16'h0000;
        rom[6][939] = 16'h0000;
        rom[6][940] = 16'h0000;
        rom[6][941] = 16'h0000;
        rom[6][942] = 16'h0000;
        rom[6][943] = 16'h0000;
        rom[6][944] = 16'h0000;
        rom[6][945] = 16'h0000;
        rom[6][946] = 16'h0000;
        rom[6][947] = 16'h0000;
        rom[6][948] = 16'h0000;
        rom[6][949] = 16'h0000;
        rom[6][950] = 16'h0000;
        rom[6][951] = 16'h0000;
        rom[6][952] = 16'h0000;
        rom[6][953] = 16'h0000;
        rom[6][954] = 16'h0000;
        rom[6][955] = 16'h0000;
        rom[6][956] = 16'h0000;
        rom[6][957] = 16'h0000;
        rom[6][958] = 16'h0000;
        rom[6][959] = 16'h0000;
        rom[6][960] = 16'h0000;
        rom[6][961] = 16'h0000;
        rom[6][962] = 16'h0000;
        rom[6][963] = 16'h0000;
        rom[6][964] = 16'h0000;
        rom[6][965] = 16'h0000;
        rom[6][966] = 16'h0000;
        rom[6][967] = 16'h0000;
        rom[6][968] = 16'h0000;
        rom[6][969] = 16'h0000;
        rom[6][970] = 16'h0000;
        rom[6][971] = 16'h0000;
        rom[6][972] = 16'h0000;
        rom[6][973] = 16'h0000;
        rom[6][974] = 16'h0000;
        rom[6][975] = 16'h0000;
        rom[6][976] = 16'h0000;
        rom[6][977] = 16'h0000;
        rom[6][978] = 16'h0000;
        rom[6][979] = 16'h0000;
        rom[6][980] = 16'hFD20;
        rom[6][981] = 16'hFD7E;
        rom[6][982] = 16'hFDC6;
        rom[6][983] = 16'hFE32;
        rom[6][984] = 16'hFE1C;
        rom[6][985] = 16'hFE15;
        rom[6][986] = 16'hFE2B;
        rom[6][987] = 16'hFEB4;
        rom[6][988] = 16'hFF27;
        rom[6][989] = 16'hFEE7;
        rom[6][990] = 16'hFEDF;
        rom[6][991] = 16'hFEF5;
        rom[6][992] = 16'hFEFC;
        rom[6][993] = 16'hFEEE;
        rom[6][994] = 16'hFF20;
        rom[6][995] = 16'hFF3D;
        rom[6][996] = 16'hFF53;
        rom[6][997] = 16'h0057;
        rom[6][998] = 16'h00EE;
        rom[6][999] = 16'h0057;
        rom[6][1000] = 16'hFFDC;
        rom[6][1001] = 16'hFFC6;
        rom[6][1002] = 16'hFF85;
        rom[6][1003] = 16'hFFEA;
        rom[6][1004] = 16'h0024;
        rom[6][1005] = 16'h0041;
        rom[6][1006] = 16'h0024;
        rom[6][1007] = 16'hFFB1;
        rom[6][1008] = 16'hFF94;
        rom[6][1009] = 16'hFE56;
        rom[6][1010] = 16'hFF53;
        rom[6][1011] = 16'hFF36;
        rom[6][1012] = 16'h0000;
        rom[6][1013] = 16'h0000;
        rom[6][1014] = 16'h0000;
        rom[6][1015] = 16'h0000;
        rom[6][1016] = 16'h0000;
        rom[6][1017] = 16'h0000;
        rom[6][1018] = 16'h0000;
        rom[6][1019] = 16'h0000;
        rom[6][1020] = 16'h0000;
        rom[6][1021] = 16'h0000;
        rom[6][1022] = 16'h0000;
        rom[6][1023] = 16'h0000;
        rom[6][1024] = 16'h0000;
        rom[6][1025] = 16'h0000;
        rom[6][1026] = 16'h0000;
        rom[6][1027] = 16'h0000;
        rom[6][1028] = 16'h0000;
        rom[6][1029] = 16'h0000;
        rom[6][1030] = 16'h0000;
        rom[6][1031] = 16'h0000;
        rom[6][1032] = 16'h0000;
        rom[6][1033] = 16'h0000;
        rom[6][1034] = 16'h0000;
        rom[6][1035] = 16'h0000;
        rom[6][1036] = 16'h0000;
        rom[6][1037] = 16'h0000;
        rom[6][1038] = 16'h0000;
        rom[6][1039] = 16'h0000;
        rom[6][1040] = 16'h0000;
        rom[6][1041] = 16'h0000;
        rom[6][1042] = 16'h0000;
        rom[6][1043] = 16'h0000;
        rom[6][1044] = 16'h0000;
        rom[6][1045] = 16'h0000;
        rom[6][1046] = 16'h0000;
        rom[6][1047] = 16'h0000;
        rom[6][1048] = 16'h0000;
        rom[6][1049] = 16'h0000;
        rom[6][1050] = 16'h0000;
        rom[6][1051] = 16'h0000;
        rom[6][1052] = 16'h0000;
        rom[6][1053] = 16'h0000;
        rom[6][1054] = 16'h0000;
        rom[6][1055] = 16'h0000;
        rom[6][1056] = 16'h0000;
        rom[6][1057] = 16'h0000;
        rom[6][1058] = 16'h0000;
        rom[6][1059] = 16'h0000;
        rom[6][1060] = 16'h0000;
        rom[6][1061] = 16'h0000;
        rom[6][1062] = 16'h0000;
        rom[6][1063] = 16'h0000;
        rom[6][1064] = 16'h0000;
        rom[6][1065] = 16'h0000;
        rom[6][1066] = 16'h0000;
        rom[6][1067] = 16'h0000;
        rom[6][1068] = 16'h0000;
        rom[6][1069] = 16'h0000;
        rom[6][1070] = 16'h0000;
        rom[6][1071] = 16'h0000;
        rom[6][1072] = 16'h0000;
        rom[6][1073] = 16'h0000;
        rom[6][1074] = 16'h0000;
        rom[6][1075] = 16'h0000;
        rom[6][1076] = 16'h0000;
        rom[6][1077] = 16'h0000;
        rom[6][1078] = 16'hFFCD;
        rom[6][1079] = 16'h0000;
        rom[6][1080] = 16'hFF9B;
        rom[6][1081] = 16'hFF53;
        rom[6][1082] = 16'hFF68;
        rom[6][1083] = 16'hFF53;
        rom[6][1084] = 16'hFE81;
        rom[6][1085] = 16'hFDA9;
        rom[6][1086] = 16'hFE15;
        rom[6][1087] = 16'hFF9B;
        rom[6][1088] = 16'h001D;
        rom[6][1089] = 16'h007B;
        rom[6][1090] = 16'h00E0;
        rom[6][1091] = 16'h0119;
        rom[6][1092] = 16'h0177;
        rom[6][1093] = 16'h0145;
        rom[6][1094] = 16'h0104;
        rom[6][1095] = 16'hFF5A;
        rom[6][1096] = 16'hFE4F;
        rom[6][1097] = 16'hFEE7;
        rom[6][1098] = 16'hFF44;
        rom[6][1099] = 16'hFF20;
        rom[6][1100] = 16'hFEA6;
        rom[6][1101] = 16'hFE41;
        rom[6][1102] = 16'hFE48;
        rom[6][1103] = 16'hFDBF;
        rom[6][1104] = 16'hFDD4;
        rom[6][1105] = 16'hFF20;
        rom[6][1106] = 16'hFFB8;
        rom[6][1107] = 16'h0016;
        rom[6][1108] = 16'hFF20;
        rom[6][1109] = 16'hFF70;
        rom[6][1110] = 16'h0000;
        rom[6][1111] = 16'h0000;
        rom[6][1112] = 16'h0000;
        rom[6][1113] = 16'h0000;
        rom[6][1114] = 16'h0000;
        rom[6][1115] = 16'h0000;
        rom[6][1116] = 16'h0000;
        rom[6][1117] = 16'h0000;
        rom[6][1118] = 16'h0000;
        rom[6][1119] = 16'h0000;
        rom[6][1120] = 16'h0000;
        rom[6][1121] = 16'h0000;
        rom[6][1122] = 16'h0000;
        rom[6][1123] = 16'h0000;
        rom[6][1124] = 16'h0000;
        rom[6][1125] = 16'h0000;
        rom[6][1126] = 16'h0000;
        rom[6][1127] = 16'h0000;
        rom[6][1128] = 16'h0000;
        rom[6][1129] = 16'h0000;
        rom[6][1130] = 16'h0000;
        rom[6][1131] = 16'h0000;
        rom[6][1132] = 16'h0000;
        rom[6][1133] = 16'h0000;
        rom[6][1134] = 16'h0000;
        rom[6][1135] = 16'h0000;
        rom[6][1136] = 16'h0000;
        rom[6][1137] = 16'h0000;
        rom[6][1138] = 16'h0000;
        rom[6][1139] = 16'h0000;
        rom[6][1140] = 16'h0000;
        rom[6][1141] = 16'h0000;
        rom[6][1142] = 16'h0000;
        rom[6][1143] = 16'h0000;
        rom[6][1144] = 16'h0000;
        rom[6][1145] = 16'h0000;
        rom[6][1146] = 16'h0000;
        rom[6][1147] = 16'h0000;
        rom[6][1148] = 16'h0000;
        rom[6][1149] = 16'h0000;
        rom[6][1150] = 16'h0000;
        rom[6][1151] = 16'h0000;
        rom[6][1152] = 16'h0000;
        rom[6][1153] = 16'h0000;
        rom[6][1154] = 16'h0000;
        rom[6][1155] = 16'h0000;
        rom[6][1156] = 16'h0000;
        rom[6][1157] = 16'h0000;
        rom[6][1158] = 16'h0000;
        rom[6][1159] = 16'h0000;
        rom[6][1160] = 16'h0000;
        rom[6][1161] = 16'h0000;
        rom[6][1162] = 16'h0000;
        rom[6][1163] = 16'h0000;
        rom[6][1164] = 16'h0000;
        rom[6][1165] = 16'h0000;
        rom[6][1166] = 16'h0000;
        rom[6][1167] = 16'h0000;
        rom[6][1168] = 16'h0000;
        rom[6][1169] = 16'h0000;
        rom[6][1170] = 16'h0000;
        rom[6][1171] = 16'h0000;
        rom[6][1172] = 16'h0000;
        rom[6][1173] = 16'h0000;
        rom[6][1174] = 16'h0000;
        rom[6][1175] = 16'h0000;
        rom[6][1176] = 16'h0313;
        rom[6][1177] = 16'hFCD0;
        rom[6][1178] = 16'hFDCD;
        rom[6][1179] = 16'hFD4B;
        rom[6][1180] = 16'hFCF5;
        rom[6][1181] = 16'hFD35;
        rom[6][1182] = 16'hFE6C;
        rom[6][1183] = 16'hFFB1;
        rom[6][1184] = 16'h00A6;
        rom[6][1185] = 16'h0048;
        rom[6][1186] = 16'hFF8D;
        rom[6][1187] = 16'hFFCD;
        rom[6][1188] = 16'hFF53;
        rom[6][1189] = 16'hFEBB;
        rom[6][1190] = 16'hFEF5;
        rom[6][1191] = 16'hFF4C;
        rom[6][1192] = 16'hFFA9;
        rom[6][1193] = 16'h0073;
        rom[6][1194] = 16'h0098;
        rom[6][1195] = 16'h0073;
        rom[6][1196] = 16'h0000;
        rom[6][1197] = 16'hFFB1;
        rom[6][1198] = 16'hFF7E;
        rom[6][1199] = 16'hFFBF;
        rom[6][1200] = 16'hFFE3;
        rom[6][1201] = 16'hFFD5;
        rom[6][1202] = 16'hFFD5;
        rom[6][1203] = 16'h0000;
        rom[6][1204] = 16'h0065;
        rom[6][1205] = 16'hFFD5;
        rom[6][1206] = 16'hFFD5;
        rom[6][1207] = 16'h003A;
        rom[6][1208] = 16'h0000;
        rom[6][1209] = 16'h0000;
        rom[6][1210] = 16'h0000;
        rom[6][1211] = 16'h0000;
        rom[6][1212] = 16'h0000;
        rom[6][1213] = 16'h0000;
        rom[6][1214] = 16'h0000;
        rom[6][1215] = 16'h0000;
        rom[6][1216] = 16'h0000;
        rom[6][1217] = 16'h0000;
        rom[6][1218] = 16'h0000;
        rom[6][1219] = 16'h0000;
        rom[6][1220] = 16'h0000;
        rom[6][1221] = 16'h0000;
        rom[6][1222] = 16'h0000;
        rom[6][1223] = 16'h0000;
        rom[6][1224] = 16'h0000;
        rom[6][1225] = 16'h0000;
        rom[6][1226] = 16'h0000;
        rom[6][1227] = 16'h0000;
        rom[6][1228] = 16'h0000;
        rom[6][1229] = 16'h0000;
        rom[6][1230] = 16'h0000;
        rom[6][1231] = 16'h0000;
        rom[6][1232] = 16'h0000;
        rom[6][1233] = 16'h0000;
        rom[6][1234] = 16'h0000;
        rom[6][1235] = 16'h0000;
        rom[6][1236] = 16'h0000;
        rom[6][1237] = 16'h0000;
        rom[6][1238] = 16'h0000;
        rom[6][1239] = 16'h0000;
        rom[6][1240] = 16'h0000;
        rom[6][1241] = 16'h0000;
        rom[6][1242] = 16'h0000;
        rom[6][1243] = 16'h0000;
        rom[6][1244] = 16'h0000;
        rom[6][1245] = 16'h0000;
        rom[6][1246] = 16'h0000;
        rom[6][1247] = 16'h0000;
        rom[6][1248] = 16'h0000;
        rom[6][1249] = 16'h0000;
        rom[6][1250] = 16'h0000;
        rom[6][1251] = 16'h0000;
        rom[6][1252] = 16'h0000;
        rom[6][1253] = 16'h0000;
        rom[6][1254] = 16'h0000;
        rom[6][1255] = 16'h0000;
        rom[6][1256] = 16'h0000;
        rom[6][1257] = 16'h0000;
        rom[6][1258] = 16'h0000;
        rom[6][1259] = 16'h0000;
        rom[6][1260] = 16'h0000;
        rom[6][1261] = 16'h0000;
        rom[6][1262] = 16'h0000;
        rom[6][1263] = 16'h0000;
        rom[6][1264] = 16'h0000;
        rom[6][1265] = 16'h0000;
        rom[6][1266] = 16'h0000;
        rom[6][1267] = 16'h0000;
        rom[6][1268] = 16'h0000;
        rom[6][1269] = 16'h0000;
        rom[6][1270] = 16'h0000;
        rom[6][1271] = 16'h0000;
        rom[6][1272] = 16'h0000;
        rom[6][1273] = 16'h0000;
        rom[7][0] = 16'h00EE;
        rom[7][1] = 16'h00F5;
        rom[7][2] = 16'h00E0;
        rom[7][3] = 16'h00AD;
        rom[7][4] = 16'h007B;
        rom[7][5] = 16'h0057;
        rom[7][6] = 16'h002B;
        rom[7][7] = 16'h000E;
        rom[7][8] = 16'hFFE3;
        rom[7][9] = 16'hFFCD;
        rom[7][10] = 16'hFFB8;
        rom[7][11] = 16'hFFA2;
        rom[7][12] = 16'hFFC6;
        rom[7][13] = 16'hFFF2;
        rom[7][14] = 16'hFFEA;
        rom[7][15] = 16'hFFD5;
        rom[7][16] = 16'h001D;
        rom[7][17] = 16'h0082;
        rom[7][18] = 16'h00B4;
        rom[7][19] = 16'h00CA;
        rom[7][20] = 16'h00D1;
        rom[7][21] = 16'h00A6;
        rom[7][22] = 16'h0090;
        rom[7][23] = 16'h00AD;
        rom[7][24] = 16'h00D9;
        rom[7][25] = 16'h00D1;
        rom[7][26] = 16'h00CA;
        rom[7][27] = 16'h012F;
        rom[7][28] = 16'h014C;
        rom[7][29] = 16'h012F;
        rom[7][30] = 16'h0104;
        rom[7][31] = 16'h0104;
        rom[7][32] = 16'h0000;
        rom[7][33] = 16'h0000;
        rom[7][34] = 16'h0000;
        rom[7][35] = 16'h0000;
        rom[7][36] = 16'h0000;
        rom[7][37] = 16'h0000;
        rom[7][38] = 16'h0000;
        rom[7][39] = 16'h0000;
        rom[7][40] = 16'h0000;
        rom[7][41] = 16'h0000;
        rom[7][42] = 16'h0000;
        rom[7][43] = 16'h0000;
        rom[7][44] = 16'h0000;
        rom[7][45] = 16'h0000;
        rom[7][46] = 16'h0000;
        rom[7][47] = 16'h0000;
        rom[7][48] = 16'h0000;
        rom[7][49] = 16'h0000;
        rom[7][50] = 16'h0000;
        rom[7][51] = 16'h0000;
        rom[7][52] = 16'h0000;
        rom[7][53] = 16'h0000;
        rom[7][54] = 16'h0000;
        rom[7][55] = 16'h0000;
        rom[7][56] = 16'h0000;
        rom[7][57] = 16'h0000;
        rom[7][58] = 16'h0000;
        rom[7][59] = 16'h0000;
        rom[7][60] = 16'h0000;
        rom[7][61] = 16'h0000;
        rom[7][62] = 16'h0000;
        rom[7][63] = 16'h0000;
        rom[7][64] = 16'h0000;
        rom[7][65] = 16'h0000;
        rom[7][66] = 16'h0000;
        rom[7][67] = 16'h0000;
        rom[7][68] = 16'h0000;
        rom[7][69] = 16'h0000;
        rom[7][70] = 16'h0000;
        rom[7][71] = 16'h0000;
        rom[7][72] = 16'h0000;
        rom[7][73] = 16'h0000;
        rom[7][74] = 16'h0000;
        rom[7][75] = 16'h0000;
        rom[7][76] = 16'h0000;
        rom[7][77] = 16'h0000;
        rom[7][78] = 16'h0000;
        rom[7][79] = 16'h0000;
        rom[7][80] = 16'h0000;
        rom[7][81] = 16'h0000;
        rom[7][82] = 16'h0000;
        rom[7][83] = 16'h0000;
        rom[7][84] = 16'h0000;
        rom[7][85] = 16'h0000;
        rom[7][86] = 16'h0000;
        rom[7][87] = 16'h0000;
        rom[7][88] = 16'h0000;
        rom[7][89] = 16'h0000;
        rom[7][90] = 16'h0000;
        rom[7][91] = 16'h0000;
        rom[7][92] = 16'h0000;
        rom[7][93] = 16'h0000;
        rom[7][94] = 16'h0000;
        rom[7][95] = 16'h0000;
        rom[7][96] = 16'h0000;
        rom[7][97] = 16'h0000;
        rom[7][98] = 16'h0200;
        rom[7][99] = 16'h0200;
        rom[7][100] = 16'h01E4;
        rom[7][101] = 16'h0186;
        rom[7][102] = 16'h0153;
        rom[7][103] = 16'h0128;
        rom[7][104] = 16'h0112;
        rom[7][105] = 16'h00F5;
        rom[7][106] = 16'h00C3;
        rom[7][107] = 16'h0098;
        rom[7][108] = 16'h0082;
        rom[7][109] = 16'h0089;
        rom[7][110] = 16'h00E7;
        rom[7][111] = 16'h010B;
        rom[7][112] = 16'h00FD;
        rom[7][113] = 16'h00CA;
        rom[7][114] = 16'h00D1;
        rom[7][115] = 16'h00C3;
        rom[7][116] = 16'h0090;
        rom[7][117] = 16'h0089;
        rom[7][118] = 16'h009F;
        rom[7][119] = 16'h0098;
        rom[7][120] = 16'hFFE3;
        rom[7][121] = 16'hFF3D;
        rom[7][122] = 16'hFF0B;
        rom[7][123] = 16'hFF61;
        rom[7][124] = 16'hFFF2;
        rom[7][125] = 16'hFF9B;
        rom[7][126] = 16'hFF9B;
        rom[7][127] = 16'h0041;
        rom[7][128] = 16'h0128;
        rom[7][129] = 16'h0186;
        rom[7][130] = 16'h0000;
        rom[7][131] = 16'h0000;
        rom[7][132] = 16'h0000;
        rom[7][133] = 16'h0000;
        rom[7][134] = 16'h0000;
        rom[7][135] = 16'h0000;
        rom[7][136] = 16'h0000;
        rom[7][137] = 16'h0000;
        rom[7][138] = 16'h0000;
        rom[7][139] = 16'h0000;
        rom[7][140] = 16'h0000;
        rom[7][141] = 16'h0000;
        rom[7][142] = 16'h0000;
        rom[7][143] = 16'h0000;
        rom[7][144] = 16'h0000;
        rom[7][145] = 16'h0000;
        rom[7][146] = 16'h0000;
        rom[7][147] = 16'h0000;
        rom[7][148] = 16'h0000;
        rom[7][149] = 16'h0000;
        rom[7][150] = 16'h0000;
        rom[7][151] = 16'h0000;
        rom[7][152] = 16'h0000;
        rom[7][153] = 16'h0000;
        rom[7][154] = 16'h0000;
        rom[7][155] = 16'h0000;
        rom[7][156] = 16'h0000;
        rom[7][157] = 16'h0000;
        rom[7][158] = 16'h0000;
        rom[7][159] = 16'h0000;
        rom[7][160] = 16'h0000;
        rom[7][161] = 16'h0000;
        rom[7][162] = 16'h0000;
        rom[7][163] = 16'h0000;
        rom[7][164] = 16'h0000;
        rom[7][165] = 16'h0000;
        rom[7][166] = 16'h0000;
        rom[7][167] = 16'h0000;
        rom[7][168] = 16'h0000;
        rom[7][169] = 16'h0000;
        rom[7][170] = 16'h0000;
        rom[7][171] = 16'h0000;
        rom[7][172] = 16'h0000;
        rom[7][173] = 16'h0000;
        rom[7][174] = 16'h0000;
        rom[7][175] = 16'h0000;
        rom[7][176] = 16'h0000;
        rom[7][177] = 16'h0000;
        rom[7][178] = 16'h0000;
        rom[7][179] = 16'h0000;
        rom[7][180] = 16'h0000;
        rom[7][181] = 16'h0000;
        rom[7][182] = 16'h0000;
        rom[7][183] = 16'h0000;
        rom[7][184] = 16'h0000;
        rom[7][185] = 16'h0000;
        rom[7][186] = 16'h0000;
        rom[7][187] = 16'h0000;
        rom[7][188] = 16'h0000;
        rom[7][189] = 16'h0000;
        rom[7][190] = 16'h0000;
        rom[7][191] = 16'h0000;
        rom[7][192] = 16'h0000;
        rom[7][193] = 16'h0000;
        rom[7][194] = 16'h0000;
        rom[7][195] = 16'h0000;
        rom[7][196] = 16'hFF94;
        rom[7][197] = 16'hFF12;
        rom[7][198] = 16'hFF2F;
        rom[7][199] = 16'hFF61;
        rom[7][200] = 16'hFF85;
        rom[7][201] = 16'hFFB1;
        rom[7][202] = 16'hFFE3;
        rom[7][203] = 16'hFFEA;
        rom[7][204] = 16'hFFEA;
        rom[7][205] = 16'h0007;
        rom[7][206] = 16'h002B;
        rom[7][207] = 16'h002B;
        rom[7][208] = 16'h0073;
        rom[7][209] = 16'h00CA;
        rom[7][210] = 16'h0112;
        rom[7][211] = 16'h0119;
        rom[7][212] = 16'h00A6;
        rom[7][213] = 16'h003A;
        rom[7][214] = 16'h0024;
        rom[7][215] = 16'h000E;
        rom[7][216] = 16'h000E;
        rom[7][217] = 16'h002B;
        rom[7][218] = 16'h0098;
        rom[7][219] = 16'h00B4;
        rom[7][220] = 16'h0089;
        rom[7][221] = 16'h0073;
        rom[7][222] = 16'h0033;
        rom[7][223] = 16'h0065;
        rom[7][224] = 16'h004F;
        rom[7][225] = 16'hFF8D;
        rom[7][226] = 16'hFECA;
        rom[7][227] = 16'hFF12;
        rom[7][228] = 16'h0000;
        rom[7][229] = 16'h0000;
        rom[7][230] = 16'h0000;
        rom[7][231] = 16'h0000;
        rom[7][232] = 16'h0000;
        rom[7][233] = 16'h0000;
        rom[7][234] = 16'h0000;
        rom[7][235] = 16'h0000;
        rom[7][236] = 16'h0000;
        rom[7][237] = 16'h0000;
        rom[7][238] = 16'h0000;
        rom[7][239] = 16'h0000;
        rom[7][240] = 16'h0000;
        rom[7][241] = 16'h0000;
        rom[7][242] = 16'h0000;
        rom[7][243] = 16'h0000;
        rom[7][244] = 16'h0000;
        rom[7][245] = 16'h0000;
        rom[7][246] = 16'h0000;
        rom[7][247] = 16'h0000;
        rom[7][248] = 16'h0000;
        rom[7][249] = 16'h0000;
        rom[7][250] = 16'h0000;
        rom[7][251] = 16'h0000;
        rom[7][252] = 16'h0000;
        rom[7][253] = 16'h0000;
        rom[7][254] = 16'h0000;
        rom[7][255] = 16'h0000;
        rom[7][256] = 16'h0000;
        rom[7][257] = 16'h0000;
        rom[7][258] = 16'h0000;
        rom[7][259] = 16'h0000;
        rom[7][260] = 16'h0000;
        rom[7][261] = 16'h0000;
        rom[7][262] = 16'h0000;
        rom[7][263] = 16'h0000;
        rom[7][264] = 16'h0000;
        rom[7][265] = 16'h0000;
        rom[7][266] = 16'h0000;
        rom[7][267] = 16'h0000;
        rom[7][268] = 16'h0000;
        rom[7][269] = 16'h0000;
        rom[7][270] = 16'h0000;
        rom[7][271] = 16'h0000;
        rom[7][272] = 16'h0000;
        rom[7][273] = 16'h0000;
        rom[7][274] = 16'h0000;
        rom[7][275] = 16'h0000;
        rom[7][276] = 16'h0000;
        rom[7][277] = 16'h0000;
        rom[7][278] = 16'h0000;
        rom[7][279] = 16'h0000;
        rom[7][280] = 16'h0000;
        rom[7][281] = 16'h0000;
        rom[7][282] = 16'h0000;
        rom[7][283] = 16'h0000;
        rom[7][284] = 16'h0000;
        rom[7][285] = 16'h0000;
        rom[7][286] = 16'h0000;
        rom[7][287] = 16'h0000;
        rom[7][288] = 16'h0000;
        rom[7][289] = 16'h0000;
        rom[7][290] = 16'h0000;
        rom[7][291] = 16'h0000;
        rom[7][292] = 16'h0000;
        rom[7][293] = 16'h0000;
        rom[7][294] = 16'h0065;
        rom[7][295] = 16'hFFF2;
        rom[7][296] = 16'hFFEA;
        rom[7][297] = 16'h002B;
        rom[7][298] = 16'h0033;
        rom[7][299] = 16'h003A;
        rom[7][300] = 16'h005E;
        rom[7][301] = 16'h0041;
        rom[7][302] = 16'h0033;
        rom[7][303] = 16'h003A;
        rom[7][304] = 16'h005E;
        rom[7][305] = 16'h0065;
        rom[7][306] = 16'h003A;
        rom[7][307] = 16'hFFB8;
        rom[7][308] = 16'hFFCD;
        rom[7][309] = 16'h003A;
        rom[7][310] = 16'hFFB1;
        rom[7][311] = 16'hFF9B;
        rom[7][312] = 16'hFF85;
        rom[7][313] = 16'hFF53;
        rom[7][314] = 16'hFF2F;
        rom[7][315] = 16'hFF12;
        rom[7][316] = 16'hFF68;
        rom[7][317] = 16'h002B;
        rom[7][318] = 16'h00AD;
        rom[7][319] = 16'h00E7;
        rom[7][320] = 16'h00A6;
        rom[7][321] = 16'h009F;
        rom[7][322] = 16'h00E0;
        rom[7][323] = 16'h0121;
        rom[7][324] = 16'h0112;
        rom[7][325] = 16'h0090;
        rom[7][326] = 16'h0000;
        rom[7][327] = 16'h0000;
        rom[7][328] = 16'h0000;
        rom[7][329] = 16'h0000;
        rom[7][330] = 16'h0000;
        rom[7][331] = 16'h0000;
        rom[7][332] = 16'h0000;
        rom[7][333] = 16'h0000;
        rom[7][334] = 16'h0000;
        rom[7][335] = 16'h0000;
        rom[7][336] = 16'h0000;
        rom[7][337] = 16'h0000;
        rom[7][338] = 16'h0000;
        rom[7][339] = 16'h0000;
        rom[7][340] = 16'h0000;
        rom[7][341] = 16'h0000;
        rom[7][342] = 16'h0000;
        rom[7][343] = 16'h0000;
        rom[7][344] = 16'h0000;
        rom[7][345] = 16'h0000;
        rom[7][346] = 16'h0000;
        rom[7][347] = 16'h0000;
        rom[7][348] = 16'h0000;
        rom[7][349] = 16'h0000;
        rom[7][350] = 16'h0000;
        rom[7][351] = 16'h0000;
        rom[7][352] = 16'h0000;
        rom[7][353] = 16'h0000;
        rom[7][354] = 16'h0000;
        rom[7][355] = 16'h0000;
        rom[7][356] = 16'h0000;
        rom[7][357] = 16'h0000;
        rom[7][358] = 16'h0000;
        rom[7][359] = 16'h0000;
        rom[7][360] = 16'h0000;
        rom[7][361] = 16'h0000;
        rom[7][362] = 16'h0000;
        rom[7][363] = 16'h0000;
        rom[7][364] = 16'h0000;
        rom[7][365] = 16'h0000;
        rom[7][366] = 16'h0000;
        rom[7][367] = 16'h0000;
        rom[7][368] = 16'h0000;
        rom[7][369] = 16'h0000;
        rom[7][370] = 16'h0000;
        rom[7][371] = 16'h0000;
        rom[7][372] = 16'h0000;
        rom[7][373] = 16'h0000;
        rom[7][374] = 16'h0000;
        rom[7][375] = 16'h0000;
        rom[7][376] = 16'h0000;
        rom[7][377] = 16'h0000;
        rom[7][378] = 16'h0000;
        rom[7][379] = 16'h0000;
        rom[7][380] = 16'h0000;
        rom[7][381] = 16'h0000;
        rom[7][382] = 16'h0000;
        rom[7][383] = 16'h0000;
        rom[7][384] = 16'h0000;
        rom[7][385] = 16'h0000;
        rom[7][386] = 16'h0000;
        rom[7][387] = 16'h0000;
        rom[7][388] = 16'h0000;
        rom[7][389] = 16'h0000;
        rom[7][390] = 16'h0000;
        rom[7][391] = 16'h0000;
        rom[7][392] = 16'h0090;
        rom[7][393] = 16'hFFF9;
        rom[7][394] = 16'hFF77;
        rom[7][395] = 16'hFFBF;
        rom[7][396] = 16'h0000;
        rom[7][397] = 16'hFFBF;
        rom[7][398] = 16'hFFB8;
        rom[7][399] = 16'h0007;
        rom[7][400] = 16'h0048;
        rom[7][401] = 16'h0065;
        rom[7][402] = 16'h0073;
        rom[7][403] = 16'h0073;
        rom[7][404] = 16'h00A6;
        rom[7][405] = 16'h00CA;
        rom[7][406] = 16'h00D1;
        rom[7][407] = 16'h00BC;
        rom[7][408] = 16'h0089;
        rom[7][409] = 16'h0073;
        rom[7][410] = 16'h0082;
        rom[7][411] = 16'h005E;
        rom[7][412] = 16'h007B;
        rom[7][413] = 16'h00B4;
        rom[7][414] = 16'h005E;
        rom[7][415] = 16'hFFD5;
        rom[7][416] = 16'hFFA2;
        rom[7][417] = 16'hFF85;
        rom[7][418] = 16'hFF20;
        rom[7][419] = 16'hFE2B;
        rom[7][420] = 16'hFE32;
        rom[7][421] = 16'hFEDF;
        rom[7][422] = 16'hFF8D;
        rom[7][423] = 16'h0033;
        rom[7][424] = 16'h0000;
        rom[7][425] = 16'h0000;
        rom[7][426] = 16'h0000;
        rom[7][427] = 16'h0000;
        rom[7][428] = 16'h0000;
        rom[7][429] = 16'h0000;
        rom[7][430] = 16'h0000;
        rom[7][431] = 16'h0000;
        rom[7][432] = 16'h0000;
        rom[7][433] = 16'h0000;
        rom[7][434] = 16'h0000;
        rom[7][435] = 16'h0000;
        rom[7][436] = 16'h0000;
        rom[7][437] = 16'h0000;
        rom[7][438] = 16'h0000;
        rom[7][439] = 16'h0000;
        rom[7][440] = 16'h0000;
        rom[7][441] = 16'h0000;
        rom[7][442] = 16'h0000;
        rom[7][443] = 16'h0000;
        rom[7][444] = 16'h0000;
        rom[7][445] = 16'h0000;
        rom[7][446] = 16'h0000;
        rom[7][447] = 16'h0000;
        rom[7][448] = 16'h0000;
        rom[7][449] = 16'h0000;
        rom[7][450] = 16'h0000;
        rom[7][451] = 16'h0000;
        rom[7][452] = 16'h0000;
        rom[7][453] = 16'h0000;
        rom[7][454] = 16'h0000;
        rom[7][455] = 16'h0000;
        rom[7][456] = 16'h0000;
        rom[7][457] = 16'h0000;
        rom[7][458] = 16'h0000;
        rom[7][459] = 16'h0000;
        rom[7][460] = 16'h0000;
        rom[7][461] = 16'h0000;
        rom[7][462] = 16'h0000;
        rom[7][463] = 16'h0000;
        rom[7][464] = 16'h0000;
        rom[7][465] = 16'h0000;
        rom[7][466] = 16'h0000;
        rom[7][467] = 16'h0000;
        rom[7][468] = 16'h0000;
        rom[7][469] = 16'h0000;
        rom[7][470] = 16'h0000;
        rom[7][471] = 16'h0000;
        rom[7][472] = 16'h0000;
        rom[7][473] = 16'h0000;
        rom[7][474] = 16'h0000;
        rom[7][475] = 16'h0000;
        rom[7][476] = 16'h0000;
        rom[7][477] = 16'h0000;
        rom[7][478] = 16'h0000;
        rom[7][479] = 16'h0000;
        rom[7][480] = 16'h0000;
        rom[7][481] = 16'h0000;
        rom[7][482] = 16'h0000;
        rom[7][483] = 16'h0000;
        rom[7][484] = 16'h0000;
        rom[7][485] = 16'h0000;
        rom[7][486] = 16'h0000;
        rom[7][487] = 16'h0000;
        rom[7][488] = 16'h0000;
        rom[7][489] = 16'h0000;
        rom[7][490] = 16'h002B;
        rom[7][491] = 16'h0065;
        rom[7][492] = 16'h0000;
        rom[7][493] = 16'h002B;
        rom[7][494] = 16'h0041;
        rom[7][495] = 16'hFFB8;
        rom[7][496] = 16'hFF68;
        rom[7][497] = 16'hFF94;
        rom[7][498] = 16'h000E;
        rom[7][499] = 16'h003A;
        rom[7][500] = 16'h0007;
        rom[7][501] = 16'h003A;
        rom[7][502] = 16'h00D1;
        rom[7][503] = 16'h00E7;
        rom[7][504] = 16'h007B;
        rom[7][505] = 16'h0016;
        rom[7][506] = 16'h007B;
        rom[7][507] = 16'h006C;
        rom[7][508] = 16'hFFF9;
        rom[7][509] = 16'hFFDC;
        rom[7][510] = 16'h0000;
        rom[7][511] = 16'h004F;
        rom[7][512] = 16'h00CA;
        rom[7][513] = 16'h005E;
        rom[7][514] = 16'h001D;
        rom[7][515] = 16'h0033;
        rom[7][516] = 16'h0065;
        rom[7][517] = 16'h009F;
        rom[7][518] = 16'h00E0;
        rom[7][519] = 16'h0121;
        rom[7][520] = 16'h0033;
        rom[7][521] = 16'hFF5A;
        rom[7][522] = 16'h0000;
        rom[7][523] = 16'h0000;
        rom[7][524] = 16'h0000;
        rom[7][525] = 16'h0000;
        rom[7][526] = 16'h0000;
        rom[7][527] = 16'h0000;
        rom[7][528] = 16'h0000;
        rom[7][529] = 16'h0000;
        rom[7][530] = 16'h0000;
        rom[7][531] = 16'h0000;
        rom[7][532] = 16'h0000;
        rom[7][533] = 16'h0000;
        rom[7][534] = 16'h0000;
        rom[7][535] = 16'h0000;
        rom[7][536] = 16'h0000;
        rom[7][537] = 16'h0000;
        rom[7][538] = 16'h0000;
        rom[7][539] = 16'h0000;
        rom[7][540] = 16'h0000;
        rom[7][541] = 16'h0000;
        rom[7][542] = 16'h0000;
        rom[7][543] = 16'h0000;
        rom[7][544] = 16'h0000;
        rom[7][545] = 16'h0000;
        rom[7][546] = 16'h0000;
        rom[7][547] = 16'h0000;
        rom[7][548] = 16'h0000;
        rom[7][549] = 16'h0000;
        rom[7][550] = 16'h0000;
        rom[7][551] = 16'h0000;
        rom[7][552] = 16'h0000;
        rom[7][553] = 16'h0000;
        rom[7][554] = 16'h0000;
        rom[7][555] = 16'h0000;
        rom[7][556] = 16'h0000;
        rom[7][557] = 16'h0000;
        rom[7][558] = 16'h0000;
        rom[7][559] = 16'h0000;
        rom[7][560] = 16'h0000;
        rom[7][561] = 16'h0000;
        rom[7][562] = 16'h0000;
        rom[7][563] = 16'h0000;
        rom[7][564] = 16'h0000;
        rom[7][565] = 16'h0000;
        rom[7][566] = 16'h0000;
        rom[7][567] = 16'h0000;
        rom[7][568] = 16'h0000;
        rom[7][569] = 16'h0000;
        rom[7][570] = 16'h0000;
        rom[7][571] = 16'h0000;
        rom[7][572] = 16'h0000;
        rom[7][573] = 16'h0000;
        rom[7][574] = 16'h0000;
        rom[7][575] = 16'h0000;
        rom[7][576] = 16'h0000;
        rom[7][577] = 16'h0000;
        rom[7][578] = 16'h0000;
        rom[7][579] = 16'h0000;
        rom[7][580] = 16'h0000;
        rom[7][581] = 16'h0000;
        rom[7][582] = 16'h0000;
        rom[7][583] = 16'h0000;
        rom[7][584] = 16'h0000;
        rom[7][585] = 16'h0000;
        rom[7][586] = 16'h0000;
        rom[7][587] = 16'h0000;
        rom[7][588] = 16'hFF19;
        rom[7][589] = 16'hFF7E;
        rom[7][590] = 16'hFF2F;
        rom[7][591] = 16'hFEFC;
        rom[7][592] = 16'hFF03;
        rom[7][593] = 16'hFEDF;
        rom[7][594] = 16'hFEE7;
        rom[7][595] = 16'hFEF5;
        rom[7][596] = 16'hFF44;
        rom[7][597] = 16'hFF70;
        rom[7][598] = 16'hFF27;
        rom[7][599] = 16'hFF61;
        rom[7][600] = 16'hFFF9;
        rom[7][601] = 16'h000E;
        rom[7][602] = 16'hFFBF;
        rom[7][603] = 16'hFF8D;
        rom[7][604] = 16'hFF61;
        rom[7][605] = 16'hFF03;
        rom[7][606] = 16'hFEF5;
        rom[7][607] = 16'hFEE7;
        rom[7][608] = 16'hFEC2;
        rom[7][609] = 16'hFF19;
        rom[7][610] = 16'hFF5A;
        rom[7][611] = 16'hFF53;
        rom[7][612] = 16'hFF27;
        rom[7][613] = 16'hFF19;
        rom[7][614] = 16'hFEBB;
        rom[7][615] = 16'hFE1C;
        rom[7][616] = 16'hFD76;
        rom[7][617] = 16'hFD3D;
        rom[7][618] = 16'hFE39;
        rom[7][619] = 16'hFEBB;
        rom[7][620] = 16'h0000;
        rom[7][621] = 16'h0000;
        rom[7][622] = 16'h0000;
        rom[7][623] = 16'h0000;
        rom[7][624] = 16'h0000;
        rom[7][625] = 16'h0000;
        rom[7][626] = 16'h0000;
        rom[7][627] = 16'h0000;
        rom[7][628] = 16'h0000;
        rom[7][629] = 16'h0000;
        rom[7][630] = 16'h0000;
        rom[7][631] = 16'h0000;
        rom[7][632] = 16'h0000;
        rom[7][633] = 16'h0000;
        rom[7][634] = 16'h0000;
        rom[7][635] = 16'h0000;
        rom[7][636] = 16'h0000;
        rom[7][637] = 16'h0000;
        rom[7][638] = 16'h0000;
        rom[7][639] = 16'h0000;
        rom[7][640] = 16'h0000;
        rom[7][641] = 16'h0000;
        rom[7][642] = 16'h0000;
        rom[7][643] = 16'h0000;
        rom[7][644] = 16'h0000;
        rom[7][645] = 16'h0000;
        rom[7][646] = 16'h0000;
        rom[7][647] = 16'h0000;
        rom[7][648] = 16'h0000;
        rom[7][649] = 16'h0000;
        rom[7][650] = 16'h0000;
        rom[7][651] = 16'h0000;
        rom[7][652] = 16'h0000;
        rom[7][653] = 16'h0000;
        rom[7][654] = 16'h0000;
        rom[7][655] = 16'h0000;
        rom[7][656] = 16'h0000;
        rom[7][657] = 16'h0000;
        rom[7][658] = 16'h0000;
        rom[7][659] = 16'h0000;
        rom[7][660] = 16'h0000;
        rom[7][661] = 16'h0000;
        rom[7][662] = 16'h0000;
        rom[7][663] = 16'h0000;
        rom[7][664] = 16'h0000;
        rom[7][665] = 16'h0000;
        rom[7][666] = 16'h0000;
        rom[7][667] = 16'h0000;
        rom[7][668] = 16'h0000;
        rom[7][669] = 16'h0000;
        rom[7][670] = 16'h0000;
        rom[7][671] = 16'h0000;
        rom[7][672] = 16'h0000;
        rom[7][673] = 16'h0000;
        rom[7][674] = 16'h0000;
        rom[7][675] = 16'h0000;
        rom[7][676] = 16'h0000;
        rom[7][677] = 16'h0000;
        rom[7][678] = 16'h0000;
        rom[7][679] = 16'h0000;
        rom[7][680] = 16'h0000;
        rom[7][681] = 16'h0000;
        rom[7][682] = 16'h0000;
        rom[7][683] = 16'h0000;
        rom[7][684] = 16'h0000;
        rom[7][685] = 16'h0000;
        rom[7][686] = 16'hFF61;
        rom[7][687] = 16'hFFCD;
        rom[7][688] = 16'hFFEA;
        rom[7][689] = 16'hFF8D;
        rom[7][690] = 16'hFF4C;
        rom[7][691] = 16'hFF8D;
        rom[7][692] = 16'hFF94;
        rom[7][693] = 16'hFFA2;
        rom[7][694] = 16'h000E;
        rom[7][695] = 16'h0033;
        rom[7][696] = 16'h0016;
        rom[7][697] = 16'h001D;
        rom[7][698] = 16'h000E;
        rom[7][699] = 16'hFFDC;
        rom[7][700] = 16'h0000;
        rom[7][701] = 16'h0048;
        rom[7][702] = 16'hFF9B;
        rom[7][703] = 16'hFFA9;
        rom[7][704] = 16'h0041;
        rom[7][705] = 16'h00B4;
        rom[7][706] = 16'h00C3;
        rom[7][707] = 16'h007B;
        rom[7][708] = 16'h0089;
        rom[7][709] = 16'h0073;
        rom[7][710] = 16'h0016;
        rom[7][711] = 16'hFF8D;
        rom[7][712] = 16'hFF5A;
        rom[7][713] = 16'hFF70;
        rom[7][714] = 16'h0007;
        rom[7][715] = 16'h005E;
        rom[7][716] = 16'h0000;
        rom[7][717] = 16'hFF53;
        rom[7][718] = 16'h0000;
        rom[7][719] = 16'h0000;
        rom[7][720] = 16'h0000;
        rom[7][721] = 16'h0000;
        rom[7][722] = 16'h0000;
        rom[7][723] = 16'h0000;
        rom[7][724] = 16'h0000;
        rom[7][725] = 16'h0000;
        rom[7][726] = 16'h0000;
        rom[7][727] = 16'h0000;
        rom[7][728] = 16'h0000;
        rom[7][729] = 16'h0000;
        rom[7][730] = 16'h0000;
        rom[7][731] = 16'h0000;
        rom[7][732] = 16'h0000;
        rom[7][733] = 16'h0000;
        rom[7][734] = 16'h0000;
        rom[7][735] = 16'h0000;
        rom[7][736] = 16'h0000;
        rom[7][737] = 16'h0000;
        rom[7][738] = 16'h0000;
        rom[7][739] = 16'h0000;
        rom[7][740] = 16'h0000;
        rom[7][741] = 16'h0000;
        rom[7][742] = 16'h0000;
        rom[7][743] = 16'h0000;
        rom[7][744] = 16'h0000;
        rom[7][745] = 16'h0000;
        rom[7][746] = 16'h0000;
        rom[7][747] = 16'h0000;
        rom[7][748] = 16'h0000;
        rom[7][749] = 16'h0000;
        rom[7][750] = 16'h0000;
        rom[7][751] = 16'h0000;
        rom[7][752] = 16'h0000;
        rom[7][753] = 16'h0000;
        rom[7][754] = 16'h0000;
        rom[7][755] = 16'h0000;
        rom[7][756] = 16'h0000;
        rom[7][757] = 16'h0000;
        rom[7][758] = 16'h0000;
        rom[7][759] = 16'h0000;
        rom[7][760] = 16'h0000;
        rom[7][761] = 16'h0000;
        rom[7][762] = 16'h0000;
        rom[7][763] = 16'h0000;
        rom[7][764] = 16'h0000;
        rom[7][765] = 16'h0000;
        rom[7][766] = 16'h0000;
        rom[7][767] = 16'h0000;
        rom[7][768] = 16'h0000;
        rom[7][769] = 16'h0000;
        rom[7][770] = 16'h0000;
        rom[7][771] = 16'h0000;
        rom[7][772] = 16'h0000;
        rom[7][773] = 16'h0000;
        rom[7][774] = 16'h0000;
        rom[7][775] = 16'h0000;
        rom[7][776] = 16'h0000;
        rom[7][777] = 16'h0000;
        rom[7][778] = 16'h0000;
        rom[7][779] = 16'h0000;
        rom[7][780] = 16'h0000;
        rom[7][781] = 16'h0000;
        rom[7][782] = 16'h0000;
        rom[7][783] = 16'h0000;
        rom[7][784] = 16'hFF61;
        rom[7][785] = 16'hFF9B;
        rom[7][786] = 16'hFF77;
        rom[7][787] = 16'hFF19;
        rom[7][788] = 16'hFEDF;
        rom[7][789] = 16'hFEF5;
        rom[7][790] = 16'hFEFC;
        rom[7][791] = 16'hFF12;
        rom[7][792] = 16'hFF5A;
        rom[7][793] = 16'hFFBF;
        rom[7][794] = 16'hFF85;
        rom[7][795] = 16'hFF7E;
        rom[7][796] = 16'hFE6C;
        rom[7][797] = 16'hFDC6;
        rom[7][798] = 16'hFDCD;
        rom[7][799] = 16'hFE6C;
        rom[7][800] = 16'hFDB0;
        rom[7][801] = 16'hFE4F;
        rom[7][802] = 16'hFFCD;
        rom[7][803] = 16'h0065;
        rom[7][804] = 16'h0073;
        rom[7][805] = 16'h0073;
        rom[7][806] = 16'h0048;
        rom[7][807] = 16'h0007;
        rom[7][808] = 16'hFFE3;
        rom[7][809] = 16'hFF61;
        rom[7][810] = 16'hFF7E;
        rom[7][811] = 16'h006C;
        rom[7][812] = 16'h00E7;
        rom[7][813] = 16'h00B4;
        rom[7][814] = 16'h00CA;
        rom[7][815] = 16'h0048;
        rom[7][816] = 16'h0000;
        rom[7][817] = 16'h0000;
        rom[7][818] = 16'h0000;
        rom[7][819] = 16'h0000;
        rom[7][820] = 16'h0000;
        rom[7][821] = 16'h0000;
        rom[7][822] = 16'h0000;
        rom[7][823] = 16'h0000;
        rom[7][824] = 16'h0000;
        rom[7][825] = 16'h0000;
        rom[7][826] = 16'h0000;
        rom[7][827] = 16'h0000;
        rom[7][828] = 16'h0000;
        rom[7][829] = 16'h0000;
        rom[7][830] = 16'h0000;
        rom[7][831] = 16'h0000;
        rom[7][832] = 16'h0000;
        rom[7][833] = 16'h0000;
        rom[7][834] = 16'h0000;
        rom[7][835] = 16'h0000;
        rom[7][836] = 16'h0000;
        rom[7][837] = 16'h0000;
        rom[7][838] = 16'h0000;
        rom[7][839] = 16'h0000;
        rom[7][840] = 16'h0000;
        rom[7][841] = 16'h0000;
        rom[7][842] = 16'h0000;
        rom[7][843] = 16'h0000;
        rom[7][844] = 16'h0000;
        rom[7][845] = 16'h0000;
        rom[7][846] = 16'h0000;
        rom[7][847] = 16'h0000;
        rom[7][848] = 16'h0000;
        rom[7][849] = 16'h0000;
        rom[7][850] = 16'h0000;
        rom[7][851] = 16'h0000;
        rom[7][852] = 16'h0000;
        rom[7][853] = 16'h0000;
        rom[7][854] = 16'h0000;
        rom[7][855] = 16'h0000;
        rom[7][856] = 16'h0000;
        rom[7][857] = 16'h0000;
        rom[7][858] = 16'h0000;
        rom[7][859] = 16'h0000;
        rom[7][860] = 16'h0000;
        rom[7][861] = 16'h0000;
        rom[7][862] = 16'h0000;
        rom[7][863] = 16'h0000;
        rom[7][864] = 16'h0000;
        rom[7][865] = 16'h0000;
        rom[7][866] = 16'h0000;
        rom[7][867] = 16'h0000;
        rom[7][868] = 16'h0000;
        rom[7][869] = 16'h0000;
        rom[7][870] = 16'h0000;
        rom[7][871] = 16'h0000;
        rom[7][872] = 16'h0000;
        rom[7][873] = 16'h0000;
        rom[7][874] = 16'h0000;
        rom[7][875] = 16'h0000;
        rom[7][876] = 16'h0000;
        rom[7][877] = 16'h0000;
        rom[7][878] = 16'h0000;
        rom[7][879] = 16'h0000;
        rom[7][880] = 16'h0000;
        rom[7][881] = 16'h0000;
        rom[7][882] = 16'hFFEA;
        rom[7][883] = 16'h012F;
        rom[7][884] = 16'h0145;
        rom[7][885] = 16'h00F5;
        rom[7][886] = 16'h0098;
        rom[7][887] = 16'h004F;
        rom[7][888] = 16'h006C;
        rom[7][889] = 16'h0082;
        rom[7][890] = 16'h0090;
        rom[7][891] = 16'h00CA;
        rom[7][892] = 16'h0090;
        rom[7][893] = 16'h004F;
        rom[7][894] = 16'hFF3D;
        rom[7][895] = 16'hFF7E;
        rom[7][896] = 16'h0024;
        rom[7][897] = 16'h006C;
        rom[7][898] = 16'h014C;
        rom[7][899] = 16'h023A;
        rom[7][900] = 16'h01B1;
        rom[7][901] = 16'h0121;
        rom[7][902] = 16'h0136;
        rom[7][903] = 16'h0153;
        rom[7][904] = 16'h00FD;
        rom[7][905] = 16'h002B;
        rom[7][906] = 16'h002B;
        rom[7][907] = 16'h002B;
        rom[7][908] = 16'h0007;
        rom[7][909] = 16'h000E;
        rom[7][910] = 16'h000E;
        rom[7][911] = 16'hFFD5;
        rom[7][912] = 16'h0016;
        rom[7][913] = 16'h001D;
        rom[7][914] = 16'h0000;
        rom[7][915] = 16'h0000;
        rom[7][916] = 16'h0000;
        rom[7][917] = 16'h0000;
        rom[7][918] = 16'h0000;
        rom[7][919] = 16'h0000;
        rom[7][920] = 16'h0000;
        rom[7][921] = 16'h0000;
        rom[7][922] = 16'h0000;
        rom[7][923] = 16'h0000;
        rom[7][924] = 16'h0000;
        rom[7][925] = 16'h0000;
        rom[7][926] = 16'h0000;
        rom[7][927] = 16'h0000;
        rom[7][928] = 16'h0000;
        rom[7][929] = 16'h0000;
        rom[7][930] = 16'h0000;
        rom[7][931] = 16'h0000;
        rom[7][932] = 16'h0000;
        rom[7][933] = 16'h0000;
        rom[7][934] = 16'h0000;
        rom[7][935] = 16'h0000;
        rom[7][936] = 16'h0000;
        rom[7][937] = 16'h0000;
        rom[7][938] = 16'h0000;
        rom[7][939] = 16'h0000;
        rom[7][940] = 16'h0000;
        rom[7][941] = 16'h0000;
        rom[7][942] = 16'h0000;
        rom[7][943] = 16'h0000;
        rom[7][944] = 16'h0000;
        rom[7][945] = 16'h0000;
        rom[7][946] = 16'h0000;
        rom[7][947] = 16'h0000;
        rom[7][948] = 16'h0000;
        rom[7][949] = 16'h0000;
        rom[7][950] = 16'h0000;
        rom[7][951] = 16'h0000;
        rom[7][952] = 16'h0000;
        rom[7][953] = 16'h0000;
        rom[7][954] = 16'h0000;
        rom[7][955] = 16'h0000;
        rom[7][956] = 16'h0000;
        rom[7][957] = 16'h0000;
        rom[7][958] = 16'h0000;
        rom[7][959] = 16'h0000;
        rom[7][960] = 16'h0000;
        rom[7][961] = 16'h0000;
        rom[7][962] = 16'h0000;
        rom[7][963] = 16'h0000;
        rom[7][964] = 16'h0000;
        rom[7][965] = 16'h0000;
        rom[7][966] = 16'h0000;
        rom[7][967] = 16'h0000;
        rom[7][968] = 16'h0000;
        rom[7][969] = 16'h0000;
        rom[7][970] = 16'h0000;
        rom[7][971] = 16'h0000;
        rom[7][972] = 16'h0000;
        rom[7][973] = 16'h0000;
        rom[7][974] = 16'h0000;
        rom[7][975] = 16'h0000;
        rom[7][976] = 16'h0000;
        rom[7][977] = 16'h0000;
        rom[7][978] = 16'h0000;
        rom[7][979] = 16'h0000;
        rom[7][980] = 16'hFF94;
        rom[7][981] = 16'hFFF9;
        rom[7][982] = 16'h001D;
        rom[7][983] = 16'h000E;
        rom[7][984] = 16'hFFE3;
        rom[7][985] = 16'hFFA9;
        rom[7][986] = 16'hFFC6;
        rom[7][987] = 16'hFFEA;
        rom[7][988] = 16'hFFEA;
        rom[7][989] = 16'hFFF9;
        rom[7][990] = 16'hFFDC;
        rom[7][991] = 16'hFFEA;
        rom[7][992] = 16'hFF4C;
        rom[7][993] = 16'hFE81;
        rom[7][994] = 16'hFDF1;
        rom[7][995] = 16'hFE0E;
        rom[7][996] = 16'hFF61;
        rom[7][997] = 16'hFFF2;
        rom[7][998] = 16'h004F;
        rom[7][999] = 16'h00A6;
        rom[7][1000] = 16'h0073;
        rom[7][1001] = 16'hFFA9;
        rom[7][1002] = 16'hFFCD;
        rom[7][1003] = 16'hFEDF;
        rom[7][1004] = 16'hFEFC;
        rom[7][1005] = 16'hFF68;
        rom[7][1006] = 16'hFF68;
        rom[7][1007] = 16'hFFA9;
        rom[7][1008] = 16'hFF2F;
        rom[7][1009] = 16'hFE89;
        rom[7][1010] = 16'hFED1;
        rom[7][1011] = 16'hFF36;
        rom[7][1012] = 16'h0000;
        rom[7][1013] = 16'h0000;
        rom[7][1014] = 16'h0000;
        rom[7][1015] = 16'h0000;
        rom[7][1016] = 16'h0000;
        rom[7][1017] = 16'h0000;
        rom[7][1018] = 16'h0000;
        rom[7][1019] = 16'h0000;
        rom[7][1020] = 16'h0000;
        rom[7][1021] = 16'h0000;
        rom[7][1022] = 16'h0000;
        rom[7][1023] = 16'h0000;
        rom[7][1024] = 16'h0000;
        rom[7][1025] = 16'h0000;
        rom[7][1026] = 16'h0000;
        rom[7][1027] = 16'h0000;
        rom[7][1028] = 16'h0000;
        rom[7][1029] = 16'h0000;
        rom[7][1030] = 16'h0000;
        rom[7][1031] = 16'h0000;
        rom[7][1032] = 16'h0000;
        rom[7][1033] = 16'h0000;
        rom[7][1034] = 16'h0000;
        rom[7][1035] = 16'h0000;
        rom[7][1036] = 16'h0000;
        rom[7][1037] = 16'h0000;
        rom[7][1038] = 16'h0000;
        rom[7][1039] = 16'h0000;
        rom[7][1040] = 16'h0000;
        rom[7][1041] = 16'h0000;
        rom[7][1042] = 16'h0000;
        rom[7][1043] = 16'h0000;
        rom[7][1044] = 16'h0000;
        rom[7][1045] = 16'h0000;
        rom[7][1046] = 16'h0000;
        rom[7][1047] = 16'h0000;
        rom[7][1048] = 16'h0000;
        rom[7][1049] = 16'h0000;
        rom[7][1050] = 16'h0000;
        rom[7][1051] = 16'h0000;
        rom[7][1052] = 16'h0000;
        rom[7][1053] = 16'h0000;
        rom[7][1054] = 16'h0000;
        rom[7][1055] = 16'h0000;
        rom[7][1056] = 16'h0000;
        rom[7][1057] = 16'h0000;
        rom[7][1058] = 16'h0000;
        rom[7][1059] = 16'h0000;
        rom[7][1060] = 16'h0000;
        rom[7][1061] = 16'h0000;
        rom[7][1062] = 16'h0000;
        rom[7][1063] = 16'h0000;
        rom[7][1064] = 16'h0000;
        rom[7][1065] = 16'h0000;
        rom[7][1066] = 16'h0000;
        rom[7][1067] = 16'h0000;
        rom[7][1068] = 16'h0000;
        rom[7][1069] = 16'h0000;
        rom[7][1070] = 16'h0000;
        rom[7][1071] = 16'h0000;
        rom[7][1072] = 16'h0000;
        rom[7][1073] = 16'h0000;
        rom[7][1074] = 16'h0000;
        rom[7][1075] = 16'h0000;
        rom[7][1076] = 16'h0000;
        rom[7][1077] = 16'h0000;
        rom[7][1078] = 16'h00EE;
        rom[7][1079] = 16'h00B4;
        rom[7][1080] = 16'h0073;
        rom[7][1081] = 16'h00A6;
        rom[7][1082] = 16'h0082;
        rom[7][1083] = 16'h0073;
        rom[7][1084] = 16'h0082;
        rom[7][1085] = 16'h0073;
        rom[7][1086] = 16'h0041;
        rom[7][1087] = 16'h002B;
        rom[7][1088] = 16'h0073;
        rom[7][1089] = 16'h0073;
        rom[7][1090] = 16'h00D1;
        rom[7][1091] = 16'h0119;
        rom[7][1092] = 16'h00CA;
        rom[7][1093] = 16'h009F;
        rom[7][1094] = 16'h00B4;
        rom[7][1095] = 16'hFFA2;
        rom[7][1096] = 16'hFF03;
        rom[7][1097] = 16'hFF3D;
        rom[7][1098] = 16'hFF44;
        rom[7][1099] = 16'hFF61;
        rom[7][1100] = 16'hFFF9;
        rom[7][1101] = 16'h005E;
        rom[7][1102] = 16'h005E;
        rom[7][1103] = 16'h0065;
        rom[7][1104] = 16'h00D9;
        rom[7][1105] = 16'h0119;
        rom[7][1106] = 16'h0162;
        rom[7][1107] = 16'h0128;
        rom[7][1108] = 16'h007B;
        rom[7][1109] = 16'hFFB1;
        rom[7][1110] = 16'h0000;
        rom[7][1111] = 16'h0000;
        rom[7][1112] = 16'h0000;
        rom[7][1113] = 16'h0000;
        rom[7][1114] = 16'h0000;
        rom[7][1115] = 16'h0000;
        rom[7][1116] = 16'h0000;
        rom[7][1117] = 16'h0000;
        rom[7][1118] = 16'h0000;
        rom[7][1119] = 16'h0000;
        rom[7][1120] = 16'h0000;
        rom[7][1121] = 16'h0000;
        rom[7][1122] = 16'h0000;
        rom[7][1123] = 16'h0000;
        rom[7][1124] = 16'h0000;
        rom[7][1125] = 16'h0000;
        rom[7][1126] = 16'h0000;
        rom[7][1127] = 16'h0000;
        rom[7][1128] = 16'h0000;
        rom[7][1129] = 16'h0000;
        rom[7][1130] = 16'h0000;
        rom[7][1131] = 16'h0000;
        rom[7][1132] = 16'h0000;
        rom[7][1133] = 16'h0000;
        rom[7][1134] = 16'h0000;
        rom[7][1135] = 16'h0000;
        rom[7][1136] = 16'h0000;
        rom[7][1137] = 16'h0000;
        rom[7][1138] = 16'h0000;
        rom[7][1139] = 16'h0000;
        rom[7][1140] = 16'h0000;
        rom[7][1141] = 16'h0000;
        rom[7][1142] = 16'h0000;
        rom[7][1143] = 16'h0000;
        rom[7][1144] = 16'h0000;
        rom[7][1145] = 16'h0000;
        rom[7][1146] = 16'h0000;
        rom[7][1147] = 16'h0000;
        rom[7][1148] = 16'h0000;
        rom[7][1149] = 16'h0000;
        rom[7][1150] = 16'h0000;
        rom[7][1151] = 16'h0000;
        rom[7][1152] = 16'h0000;
        rom[7][1153] = 16'h0000;
        rom[7][1154] = 16'h0000;
        rom[7][1155] = 16'h0000;
        rom[7][1156] = 16'h0000;
        rom[7][1157] = 16'h0000;
        rom[7][1158] = 16'h0000;
        rom[7][1159] = 16'h0000;
        rom[7][1160] = 16'h0000;
        rom[7][1161] = 16'h0000;
        rom[7][1162] = 16'h0000;
        rom[7][1163] = 16'h0000;
        rom[7][1164] = 16'h0000;
        rom[7][1165] = 16'h0000;
        rom[7][1166] = 16'h0000;
        rom[7][1167] = 16'h0000;
        rom[7][1168] = 16'h0000;
        rom[7][1169] = 16'h0000;
        rom[7][1170] = 16'h0000;
        rom[7][1171] = 16'h0000;
        rom[7][1172] = 16'h0000;
        rom[7][1173] = 16'h0000;
        rom[7][1174] = 16'h0000;
        rom[7][1175] = 16'h0000;
        rom[7][1176] = 16'h0112;
        rom[7][1177] = 16'h003A;
        rom[7][1178] = 16'hFFF2;
        rom[7][1179] = 16'hFF85;
        rom[7][1180] = 16'hFF4C;
        rom[7][1181] = 16'hFF20;
        rom[7][1182] = 16'hFFB1;
        rom[7][1183] = 16'h000E;
        rom[7][1184] = 16'hFFC6;
        rom[7][1185] = 16'hFF85;
        rom[7][1186] = 16'hFFA9;
        rom[7][1187] = 16'hFFD5;
        rom[7][1188] = 16'hFF8D;
        rom[7][1189] = 16'hFE41;
        rom[7][1190] = 16'hFD9B;
        rom[7][1191] = 16'hFE2B;
        rom[7][1192] = 16'hFE32;
        rom[7][1193] = 16'hFE89;
        rom[7][1194] = 16'hFE65;
        rom[7][1195] = 16'hFE81;
        rom[7][1196] = 16'hFE97;
        rom[7][1197] = 16'hFE97;
        rom[7][1198] = 16'hFF19;
        rom[7][1199] = 16'hFF85;
        rom[7][1200] = 16'hFF94;
        rom[7][1201] = 16'hFFBF;
        rom[7][1202] = 16'hFF70;
        rom[7][1203] = 16'hFF2F;
        rom[7][1204] = 16'hFEFC;
        rom[7][1205] = 16'hFE73;
        rom[7][1206] = 16'hFF27;
        rom[7][1207] = 16'hFFBF;
        rom[7][1208] = 16'h0000;
        rom[7][1209] = 16'h0000;
        rom[7][1210] = 16'h0000;
        rom[7][1211] = 16'h0000;
        rom[7][1212] = 16'h0000;
        rom[7][1213] = 16'h0000;
        rom[7][1214] = 16'h0000;
        rom[7][1215] = 16'h0000;
        rom[7][1216] = 16'h0000;
        rom[7][1217] = 16'h0000;
        rom[7][1218] = 16'h0000;
        rom[7][1219] = 16'h0000;
        rom[7][1220] = 16'h0000;
        rom[7][1221] = 16'h0000;
        rom[7][1222] = 16'h0000;
        rom[7][1223] = 16'h0000;
        rom[7][1224] = 16'h0000;
        rom[7][1225] = 16'h0000;
        rom[7][1226] = 16'h0000;
        rom[7][1227] = 16'h0000;
        rom[7][1228] = 16'h0000;
        rom[7][1229] = 16'h0000;
        rom[7][1230] = 16'h0000;
        rom[7][1231] = 16'h0000;
        rom[7][1232] = 16'h0000;
        rom[7][1233] = 16'h0000;
        rom[7][1234] = 16'h0000;
        rom[7][1235] = 16'h0000;
        rom[7][1236] = 16'h0000;
        rom[7][1237] = 16'h0000;
        rom[7][1238] = 16'h0000;
        rom[7][1239] = 16'h0000;
        rom[7][1240] = 16'h0000;
        rom[7][1241] = 16'h0000;
        rom[7][1242] = 16'h0000;
        rom[7][1243] = 16'h0000;
        rom[7][1244] = 16'h0000;
        rom[7][1245] = 16'h0000;
        rom[7][1246] = 16'h0000;
        rom[7][1247] = 16'h0000;
        rom[7][1248] = 16'h0000;
        rom[7][1249] = 16'h0000;
        rom[7][1250] = 16'h0000;
        rom[7][1251] = 16'h0000;
        rom[7][1252] = 16'h0000;
        rom[7][1253] = 16'h0000;
        rom[7][1254] = 16'h0000;
        rom[7][1255] = 16'h0000;
        rom[7][1256] = 16'h0000;
        rom[7][1257] = 16'h0000;
        rom[7][1258] = 16'h0000;
        rom[7][1259] = 16'h0000;
        rom[7][1260] = 16'h0000;
        rom[7][1261] = 16'h0000;
        rom[7][1262] = 16'h0000;
        rom[7][1263] = 16'h0000;
        rom[7][1264] = 16'h0000;
        rom[7][1265] = 16'h0000;
        rom[7][1266] = 16'h0000;
        rom[7][1267] = 16'h0000;
        rom[7][1268] = 16'h0000;
        rom[7][1269] = 16'h0000;
        rom[7][1270] = 16'h0000;
        rom[7][1271] = 16'h0000;
        rom[7][1272] = 16'h0000;
        rom[7][1273] = 16'h0000;
        rom[8][0] = 16'hFF68;
        rom[8][1] = 16'hFF77;
        rom[8][2] = 16'hFF77;
        rom[8][3] = 16'hFFBF;
        rom[8][4] = 16'hFFF9;
        rom[8][5] = 16'hFFF9;
        rom[8][6] = 16'hFFDC;
        rom[8][7] = 16'hFFB1;
        rom[8][8] = 16'hFF5A;
        rom[8][9] = 16'hFF8D;
        rom[8][10] = 16'h0000;
        rom[8][11] = 16'h0024;
        rom[8][12] = 16'h0007;
        rom[8][13] = 16'hFFE3;
        rom[8][14] = 16'hFFD5;
        rom[8][15] = 16'hFFEA;
        rom[8][16] = 16'hFFCD;
        rom[8][17] = 16'hFF70;
        rom[8][18] = 16'hFEF5;
        rom[8][19] = 16'hFF68;
        rom[8][20] = 16'hFFA2;
        rom[8][21] = 16'hFF68;
        rom[8][22] = 16'hFF19;
        rom[8][23] = 16'hFEEE;
        rom[8][24] = 16'hFEFC;
        rom[8][25] = 16'hFF0B;
        rom[8][26] = 16'hFF20;
        rom[8][27] = 16'hFF27;
        rom[8][28] = 16'hFF3D;
        rom[8][29] = 16'hFF44;
        rom[8][30] = 16'hFF5A;
        rom[8][31] = 16'hFF4C;
        rom[8][32] = 16'h0000;
        rom[8][33] = 16'h0000;
        rom[8][34] = 16'h0000;
        rom[8][35] = 16'h0000;
        rom[8][36] = 16'h0000;
        rom[8][37] = 16'h0000;
        rom[8][38] = 16'h0000;
        rom[8][39] = 16'h0000;
        rom[8][40] = 16'h0000;
        rom[8][41] = 16'h0000;
        rom[8][42] = 16'h0000;
        rom[8][43] = 16'h0000;
        rom[8][44] = 16'h0000;
        rom[8][45] = 16'h0000;
        rom[8][46] = 16'h0000;
        rom[8][47] = 16'h0000;
        rom[8][48] = 16'h0000;
        rom[8][49] = 16'h0000;
        rom[8][50] = 16'h0000;
        rom[8][51] = 16'h0000;
        rom[8][52] = 16'h0000;
        rom[8][53] = 16'h0000;
        rom[8][54] = 16'h0000;
        rom[8][55] = 16'h0000;
        rom[8][56] = 16'h0000;
        rom[8][57] = 16'h0000;
        rom[8][58] = 16'h0000;
        rom[8][59] = 16'h0000;
        rom[8][60] = 16'h0000;
        rom[8][61] = 16'h0000;
        rom[8][62] = 16'h0000;
        rom[8][63] = 16'h0000;
        rom[8][64] = 16'h0000;
        rom[8][65] = 16'h0000;
        rom[8][66] = 16'h0000;
        rom[8][67] = 16'h0000;
        rom[8][68] = 16'h0000;
        rom[8][69] = 16'h0000;
        rom[8][70] = 16'h0000;
        rom[8][71] = 16'h0000;
        rom[8][72] = 16'h0000;
        rom[8][73] = 16'h0000;
        rom[8][74] = 16'h0000;
        rom[8][75] = 16'h0000;
        rom[8][76] = 16'h0000;
        rom[8][77] = 16'h0000;
        rom[8][78] = 16'h0000;
        rom[8][79] = 16'h0000;
        rom[8][80] = 16'h0000;
        rom[8][81] = 16'h0000;
        rom[8][82] = 16'h0000;
        rom[8][83] = 16'h0000;
        rom[8][84] = 16'h0000;
        rom[8][85] = 16'h0000;
        rom[8][86] = 16'h0000;
        rom[8][87] = 16'h0000;
        rom[8][88] = 16'h0000;
        rom[8][89] = 16'h0000;
        rom[8][90] = 16'h0000;
        rom[8][91] = 16'h0000;
        rom[8][92] = 16'h0000;
        rom[8][93] = 16'h0000;
        rom[8][94] = 16'h0000;
        rom[8][95] = 16'h0000;
        rom[8][96] = 16'h0000;
        rom[8][97] = 16'h0000;
        rom[8][98] = 16'h018D;
        rom[8][99] = 16'h0194;
        rom[8][100] = 16'h017F;
        rom[8][101] = 16'h012F;
        rom[8][102] = 16'h0112;
        rom[8][103] = 16'h00D1;
        rom[8][104] = 16'h0090;
        rom[8][105] = 16'h0065;
        rom[8][106] = 16'h003A;
        rom[8][107] = 16'h0162;
        rom[8][108] = 16'h0208;
        rom[8][109] = 16'h0225;
        rom[8][110] = 16'h01F9;
        rom[8][111] = 16'h01C7;
        rom[8][112] = 16'h01BF;
        rom[8][113] = 16'h01EB;
        rom[8][114] = 16'h01DC;
        rom[8][115] = 16'h0194;
        rom[8][116] = 16'h0104;
        rom[8][117] = 16'h0119;
        rom[8][118] = 16'h0136;
        rom[8][119] = 16'h00EE;
        rom[8][120] = 16'h00B4;
        rom[8][121] = 16'h007B;
        rom[8][122] = 16'h006C;
        rom[8][123] = 16'h007B;
        rom[8][124] = 16'h007B;
        rom[8][125] = 16'h0082;
        rom[8][126] = 16'h009F;
        rom[8][127] = 16'h0098;
        rom[8][128] = 16'h00BC;
        rom[8][129] = 16'h00B4;
        rom[8][130] = 16'h0000;
        rom[8][131] = 16'h0000;
        rom[8][132] = 16'h0000;
        rom[8][133] = 16'h0000;
        rom[8][134] = 16'h0000;
        rom[8][135] = 16'h0000;
        rom[8][136] = 16'h0000;
        rom[8][137] = 16'h0000;
        rom[8][138] = 16'h0000;
        rom[8][139] = 16'h0000;
        rom[8][140] = 16'h0000;
        rom[8][141] = 16'h0000;
        rom[8][142] = 16'h0000;
        rom[8][143] = 16'h0000;
        rom[8][144] = 16'h0000;
        rom[8][145] = 16'h0000;
        rom[8][146] = 16'h0000;
        rom[8][147] = 16'h0000;
        rom[8][148] = 16'h0000;
        rom[8][149] = 16'h0000;
        rom[8][150] = 16'h0000;
        rom[8][151] = 16'h0000;
        rom[8][152] = 16'h0000;
        rom[8][153] = 16'h0000;
        rom[8][154] = 16'h0000;
        rom[8][155] = 16'h0000;
        rom[8][156] = 16'h0000;
        rom[8][157] = 16'h0000;
        rom[8][158] = 16'h0000;
        rom[8][159] = 16'h0000;
        rom[8][160] = 16'h0000;
        rom[8][161] = 16'h0000;
        rom[8][162] = 16'h0000;
        rom[8][163] = 16'h0000;
        rom[8][164] = 16'h0000;
        rom[8][165] = 16'h0000;
        rom[8][166] = 16'h0000;
        rom[8][167] = 16'h0000;
        rom[8][168] = 16'h0000;
        rom[8][169] = 16'h0000;
        rom[8][170] = 16'h0000;
        rom[8][171] = 16'h0000;
        rom[8][172] = 16'h0000;
        rom[8][173] = 16'h0000;
        rom[8][174] = 16'h0000;
        rom[8][175] = 16'h0000;
        rom[8][176] = 16'h0000;
        rom[8][177] = 16'h0000;
        rom[8][178] = 16'h0000;
        rom[8][179] = 16'h0000;
        rom[8][180] = 16'h0000;
        rom[8][181] = 16'h0000;
        rom[8][182] = 16'h0000;
        rom[8][183] = 16'h0000;
        rom[8][184] = 16'h0000;
        rom[8][185] = 16'h0000;
        rom[8][186] = 16'h0000;
        rom[8][187] = 16'h0000;
        rom[8][188] = 16'h0000;
        rom[8][189] = 16'h0000;
        rom[8][190] = 16'h0000;
        rom[8][191] = 16'h0000;
        rom[8][192] = 16'h0000;
        rom[8][193] = 16'h0000;
        rom[8][194] = 16'h0000;
        rom[8][195] = 16'h0000;
        rom[8][196] = 16'h0000;
        rom[8][197] = 16'hFFA2;
        rom[8][198] = 16'hFF7E;
        rom[8][199] = 16'hFE65;
        rom[8][200] = 16'hFDA2;
        rom[8][201] = 16'hFD6F;
        rom[8][202] = 16'hFD52;
        rom[8][203] = 16'hFDA9;
        rom[8][204] = 16'hFE73;
        rom[8][205] = 16'hFF5A;
        rom[8][206] = 16'hFEE7;
        rom[8][207] = 16'hFE7A;
        rom[8][208] = 16'hFE4F;
        rom[8][209] = 16'hFE56;
        rom[8][210] = 16'hFE5D;
        rom[8][211] = 16'hFE6C;
        rom[8][212] = 16'hFEA6;
        rom[8][213] = 16'hFF27;
        rom[8][214] = 16'hFF61;
        rom[8][215] = 16'hFECA;
        rom[8][216] = 16'hFE81;
        rom[8][217] = 16'hFEB4;
        rom[8][218] = 16'hFF36;
        rom[8][219] = 16'hFF5A;
        rom[8][220] = 16'hFF3D;
        rom[8][221] = 16'hFF3D;
        rom[8][222] = 16'hFF12;
        rom[8][223] = 16'hFF03;
        rom[8][224] = 16'hFF19;
        rom[8][225] = 16'hFEC2;
        rom[8][226] = 16'hFE90;
        rom[8][227] = 16'hFE9E;
        rom[8][228] = 16'h0000;
        rom[8][229] = 16'h0000;
        rom[8][230] = 16'h0000;
        rom[8][231] = 16'h0000;
        rom[8][232] = 16'h0000;
        rom[8][233] = 16'h0000;
        rom[8][234] = 16'h0000;
        rom[8][235] = 16'h0000;
        rom[8][236] = 16'h0000;
        rom[8][237] = 16'h0000;
        rom[8][238] = 16'h0000;
        rom[8][239] = 16'h0000;
        rom[8][240] = 16'h0000;
        rom[8][241] = 16'h0000;
        rom[8][242] = 16'h0000;
        rom[8][243] = 16'h0000;
        rom[8][244] = 16'h0000;
        rom[8][245] = 16'h0000;
        rom[8][246] = 16'h0000;
        rom[8][247] = 16'h0000;
        rom[8][248] = 16'h0000;
        rom[8][249] = 16'h0000;
        rom[8][250] = 16'h0000;
        rom[8][251] = 16'h0000;
        rom[8][252] = 16'h0000;
        rom[8][253] = 16'h0000;
        rom[8][254] = 16'h0000;
        rom[8][255] = 16'h0000;
        rom[8][256] = 16'h0000;
        rom[8][257] = 16'h0000;
        rom[8][258] = 16'h0000;
        rom[8][259] = 16'h0000;
        rom[8][260] = 16'h0000;
        rom[8][261] = 16'h0000;
        rom[8][262] = 16'h0000;
        rom[8][263] = 16'h0000;
        rom[8][264] = 16'h0000;
        rom[8][265] = 16'h0000;
        rom[8][266] = 16'h0000;
        rom[8][267] = 16'h0000;
        rom[8][268] = 16'h0000;
        rom[8][269] = 16'h0000;
        rom[8][270] = 16'h0000;
        rom[8][271] = 16'h0000;
        rom[8][272] = 16'h0000;
        rom[8][273] = 16'h0000;
        rom[8][274] = 16'h0000;
        rom[8][275] = 16'h0000;
        rom[8][276] = 16'h0000;
        rom[8][277] = 16'h0000;
        rom[8][278] = 16'h0000;
        rom[8][279] = 16'h0000;
        rom[8][280] = 16'h0000;
        rom[8][281] = 16'h0000;
        rom[8][282] = 16'h0000;
        rom[8][283] = 16'h0000;
        rom[8][284] = 16'h0000;
        rom[8][285] = 16'h0000;
        rom[8][286] = 16'h0000;
        rom[8][287] = 16'h0000;
        rom[8][288] = 16'h0000;
        rom[8][289] = 16'h0000;
        rom[8][290] = 16'h0000;
        rom[8][291] = 16'h0000;
        rom[8][292] = 16'h0000;
        rom[8][293] = 16'h0000;
        rom[8][294] = 16'hFEEE;
        rom[8][295] = 16'hFF27;
        rom[8][296] = 16'hFF4C;
        rom[8][297] = 16'hFFCD;
        rom[8][298] = 16'h000E;
        rom[8][299] = 16'h005E;
        rom[8][300] = 16'h007B;
        rom[8][301] = 16'h009F;
        rom[8][302] = 16'h00D1;
        rom[8][303] = 16'hFFDC;
        rom[8][304] = 16'hFFEA;
        rom[8][305] = 16'hFFC6;
        rom[8][306] = 16'hFF68;
        rom[8][307] = 16'hFF27;
        rom[8][308] = 16'hFF0B;
        rom[8][309] = 16'hFF0B;
        rom[8][310] = 16'hFF3D;
        rom[8][311] = 16'hFF44;
        rom[8][312] = 16'hFF20;
        rom[8][313] = 16'hFFC6;
        rom[8][314] = 16'h000E;
        rom[8][315] = 16'hFFDC;
        rom[8][316] = 16'hFF94;
        rom[8][317] = 16'hFFB1;
        rom[8][318] = 16'hFFF9;
        rom[8][319] = 16'hFFF9;
        rom[8][320] = 16'hFFB8;
        rom[8][321] = 16'hFFB8;
        rom[8][322] = 16'hFFDC;
        rom[8][323] = 16'hFF9B;
        rom[8][324] = 16'hFF3D;
        rom[8][325] = 16'hFF2F;
        rom[8][326] = 16'h0000;
        rom[8][327] = 16'h0000;
        rom[8][328] = 16'h0000;
        rom[8][329] = 16'h0000;
        rom[8][330] = 16'h0000;
        rom[8][331] = 16'h0000;
        rom[8][332] = 16'h0000;
        rom[8][333] = 16'h0000;
        rom[8][334] = 16'h0000;
        rom[8][335] = 16'h0000;
        rom[8][336] = 16'h0000;
        rom[8][337] = 16'h0000;
        rom[8][338] = 16'h0000;
        rom[8][339] = 16'h0000;
        rom[8][340] = 16'h0000;
        rom[8][341] = 16'h0000;
        rom[8][342] = 16'h0000;
        rom[8][343] = 16'h0000;
        rom[8][344] = 16'h0000;
        rom[8][345] = 16'h0000;
        rom[8][346] = 16'h0000;
        rom[8][347] = 16'h0000;
        rom[8][348] = 16'h0000;
        rom[8][349] = 16'h0000;
        rom[8][350] = 16'h0000;
        rom[8][351] = 16'h0000;
        rom[8][352] = 16'h0000;
        rom[8][353] = 16'h0000;
        rom[8][354] = 16'h0000;
        rom[8][355] = 16'h0000;
        rom[8][356] = 16'h0000;
        rom[8][357] = 16'h0000;
        rom[8][358] = 16'h0000;
        rom[8][359] = 16'h0000;
        rom[8][360] = 16'h0000;
        rom[8][361] = 16'h0000;
        rom[8][362] = 16'h0000;
        rom[8][363] = 16'h0000;
        rom[8][364] = 16'h0000;
        rom[8][365] = 16'h0000;
        rom[8][366] = 16'h0000;
        rom[8][367] = 16'h0000;
        rom[8][368] = 16'h0000;
        rom[8][369] = 16'h0000;
        rom[8][370] = 16'h0000;
        rom[8][371] = 16'h0000;
        rom[8][372] = 16'h0000;
        rom[8][373] = 16'h0000;
        rom[8][374] = 16'h0000;
        rom[8][375] = 16'h0000;
        rom[8][376] = 16'h0000;
        rom[8][377] = 16'h0000;
        rom[8][378] = 16'h0000;
        rom[8][379] = 16'h0000;
        rom[8][380] = 16'h0000;
        rom[8][381] = 16'h0000;
        rom[8][382] = 16'h0000;
        rom[8][383] = 16'h0000;
        rom[8][384] = 16'h0000;
        rom[8][385] = 16'h0000;
        rom[8][386] = 16'h0000;
        rom[8][387] = 16'h0000;
        rom[8][388] = 16'h0000;
        rom[8][389] = 16'h0000;
        rom[8][390] = 16'h0000;
        rom[8][391] = 16'h0000;
        rom[8][392] = 16'hFF0B;
        rom[8][393] = 16'hFF53;
        rom[8][394] = 16'hFF7E;
        rom[8][395] = 16'hFE89;
        rom[8][396] = 16'hFE0E;
        rom[8][397] = 16'hFE07;
        rom[8][398] = 16'hFE4F;
        rom[8][399] = 16'hFEDF;
        rom[8][400] = 16'hFFB8;
        rom[8][401] = 16'hFF7E;
        rom[8][402] = 16'hFF27;
        rom[8][403] = 16'hFEFC;
        rom[8][404] = 16'hFEF5;
        rom[8][405] = 16'hFEFC;
        rom[8][406] = 16'hFEDF;
        rom[8][407] = 16'hFEAD;
        rom[8][408] = 16'hFEC2;
        rom[8][409] = 16'hFF0B;
        rom[8][410] = 16'hFF9B;
        rom[8][411] = 16'hFEA6;
        rom[8][412] = 16'hFEA6;
        rom[8][413] = 16'hFEFC;
        rom[8][414] = 16'hFF5A;
        rom[8][415] = 16'h0000;
        rom[8][416] = 16'h0082;
        rom[8][417] = 16'h0090;
        rom[8][418] = 16'h003A;
        rom[8][419] = 16'h000E;
        rom[8][420] = 16'h0033;
        rom[8][421] = 16'h003A;
        rom[8][422] = 16'hFFF2;
        rom[8][423] = 16'h000E;
        rom[8][424] = 16'h0000;
        rom[8][425] = 16'h0000;
        rom[8][426] = 16'h0000;
        rom[8][427] = 16'h0000;
        rom[8][428] = 16'h0000;
        rom[8][429] = 16'h0000;
        rom[8][430] = 16'h0000;
        rom[8][431] = 16'h0000;
        rom[8][432] = 16'h0000;
        rom[8][433] = 16'h0000;
        rom[8][434] = 16'h0000;
        rom[8][435] = 16'h0000;
        rom[8][436] = 16'h0000;
        rom[8][437] = 16'h0000;
        rom[8][438] = 16'h0000;
        rom[8][439] = 16'h0000;
        rom[8][440] = 16'h0000;
        rom[8][441] = 16'h0000;
        rom[8][442] = 16'h0000;
        rom[8][443] = 16'h0000;
        rom[8][444] = 16'h0000;
        rom[8][445] = 16'h0000;
        rom[8][446] = 16'h0000;
        rom[8][447] = 16'h0000;
        rom[8][448] = 16'h0000;
        rom[8][449] = 16'h0000;
        rom[8][450] = 16'h0000;
        rom[8][451] = 16'h0000;
        rom[8][452] = 16'h0000;
        rom[8][453] = 16'h0000;
        rom[8][454] = 16'h0000;
        rom[8][455] = 16'h0000;
        rom[8][456] = 16'h0000;
        rom[8][457] = 16'h0000;
        rom[8][458] = 16'h0000;
        rom[8][459] = 16'h0000;
        rom[8][460] = 16'h0000;
        rom[8][461] = 16'h0000;
        rom[8][462] = 16'h0000;
        rom[8][463] = 16'h0000;
        rom[8][464] = 16'h0000;
        rom[8][465] = 16'h0000;
        rom[8][466] = 16'h0000;
        rom[8][467] = 16'h0000;
        rom[8][468] = 16'h0000;
        rom[8][469] = 16'h0000;
        rom[8][470] = 16'h0000;
        rom[8][471] = 16'h0000;
        rom[8][472] = 16'h0000;
        rom[8][473] = 16'h0000;
        rom[8][474] = 16'h0000;
        rom[8][475] = 16'h0000;
        rom[8][476] = 16'h0000;
        rom[8][477] = 16'h0000;
        rom[8][478] = 16'h0000;
        rom[8][479] = 16'h0000;
        rom[8][480] = 16'h0000;
        rom[8][481] = 16'h0000;
        rom[8][482] = 16'h0000;
        rom[8][483] = 16'h0000;
        rom[8][484] = 16'h0000;
        rom[8][485] = 16'h0000;
        rom[8][486] = 16'h0000;
        rom[8][487] = 16'h0000;
        rom[8][488] = 16'h0000;
        rom[8][489] = 16'h0000;
        rom[8][490] = 16'hFE4F;
        rom[8][491] = 16'hFE48;
        rom[8][492] = 16'hFE4F;
        rom[8][493] = 16'hFE15;
        rom[8][494] = 16'hFDB0;
        rom[8][495] = 16'hFD61;
        rom[8][496] = 16'hFD4B;
        rom[8][497] = 16'hFDB0;
        rom[8][498] = 16'hFE4F;
        rom[8][499] = 16'hFE48;
        rom[8][500] = 16'hFDF8;
        rom[8][501] = 16'hFE07;
        rom[8][502] = 16'hFE65;
        rom[8][503] = 16'hFED8;
        rom[8][504] = 16'hFEEE;
        rom[8][505] = 16'hFEC2;
        rom[8][506] = 16'hFEA6;
        rom[8][507] = 16'hFECA;
        rom[8][508] = 16'hFF19;
        rom[8][509] = 16'hFDB7;
        rom[8][510] = 16'hFD6F;
        rom[8][511] = 16'hFD8C;
        rom[8][512] = 16'hFDEA;
        rom[8][513] = 16'hFE73;
        rom[8][514] = 16'hFEE7;
        rom[8][515] = 16'hFF27;
        rom[8][516] = 16'hFEE7;
        rom[8][517] = 16'hFEB4;
        rom[8][518] = 16'hFED8;
        rom[8][519] = 16'hFF0B;
        rom[8][520] = 16'hFEA6;
        rom[8][521] = 16'hFEBB;
        rom[8][522] = 16'h0000;
        rom[8][523] = 16'h0000;
        rom[8][524] = 16'h0000;
        rom[8][525] = 16'h0000;
        rom[8][526] = 16'h0000;
        rom[8][527] = 16'h0000;
        rom[8][528] = 16'h0000;
        rom[8][529] = 16'h0000;
        rom[8][530] = 16'h0000;
        rom[8][531] = 16'h0000;
        rom[8][532] = 16'h0000;
        rom[8][533] = 16'h0000;
        rom[8][534] = 16'h0000;
        rom[8][535] = 16'h0000;
        rom[8][536] = 16'h0000;
        rom[8][537] = 16'h0000;
        rom[8][538] = 16'h0000;
        rom[8][539] = 16'h0000;
        rom[8][540] = 16'h0000;
        rom[8][541] = 16'h0000;
        rom[8][542] = 16'h0000;
        rom[8][543] = 16'h0000;
        rom[8][544] = 16'h0000;
        rom[8][545] = 16'h0000;
        rom[8][546] = 16'h0000;
        rom[8][547] = 16'h0000;
        rom[8][548] = 16'h0000;
        rom[8][549] = 16'h0000;
        rom[8][550] = 16'h0000;
        rom[8][551] = 16'h0000;
        rom[8][552] = 16'h0000;
        rom[8][553] = 16'h0000;
        rom[8][554] = 16'h0000;
        rom[8][555] = 16'h0000;
        rom[8][556] = 16'h0000;
        rom[8][557] = 16'h0000;
        rom[8][558] = 16'h0000;
        rom[8][559] = 16'h0000;
        rom[8][560] = 16'h0000;
        rom[8][561] = 16'h0000;
        rom[8][562] = 16'h0000;
        rom[8][563] = 16'h0000;
        rom[8][564] = 16'h0000;
        rom[8][565] = 16'h0000;
        rom[8][566] = 16'h0000;
        rom[8][567] = 16'h0000;
        rom[8][568] = 16'h0000;
        rom[8][569] = 16'h0000;
        rom[8][570] = 16'h0000;
        rom[8][571] = 16'h0000;
        rom[8][572] = 16'h0000;
        rom[8][573] = 16'h0000;
        rom[8][574] = 16'h0000;
        rom[8][575] = 16'h0000;
        rom[8][576] = 16'h0000;
        rom[8][577] = 16'h0000;
        rom[8][578] = 16'h0000;
        rom[8][579] = 16'h0000;
        rom[8][580] = 16'h0000;
        rom[8][581] = 16'h0000;
        rom[8][582] = 16'h0000;
        rom[8][583] = 16'h0000;
        rom[8][584] = 16'h0000;
        rom[8][585] = 16'h0000;
        rom[8][586] = 16'h0000;
        rom[8][587] = 16'h0000;
        rom[8][588] = 16'hFF19;
        rom[8][589] = 16'hFF9B;
        rom[8][590] = 16'hFFDC;
        rom[8][591] = 16'h0170;
        rom[8][592] = 16'h0233;
        rom[8][593] = 16'h0208;
        rom[8][594] = 16'h0225;
        rom[8][595] = 16'h0233;
        rom[8][596] = 16'h0194;
        rom[8][597] = 16'h00CA;
        rom[8][598] = 16'h0128;
        rom[8][599] = 16'h0177;
        rom[8][600] = 16'h01D5;
        rom[8][601] = 16'h0233;
        rom[8][602] = 16'h0250;
        rom[8][603] = 16'h0257;
        rom[8][604] = 16'h021D;
        rom[8][605] = 16'h01B1;
        rom[8][606] = 16'h0162;
        rom[8][607] = 16'h0170;
        rom[8][608] = 16'h015A;
        rom[8][609] = 16'h00E7;
        rom[8][610] = 16'h0057;
        rom[8][611] = 16'h0024;
        rom[8][612] = 16'h004F;
        rom[8][613] = 16'h0065;
        rom[8][614] = 16'h005E;
        rom[8][615] = 16'h0082;
        rom[8][616] = 16'h009F;
        rom[8][617] = 16'h00C3;
        rom[8][618] = 16'h0057;
        rom[8][619] = 16'hFFBF;
        rom[8][620] = 16'h0000;
        rom[8][621] = 16'h0000;
        rom[8][622] = 16'h0000;
        rom[8][623] = 16'h0000;
        rom[8][624] = 16'h0000;
        rom[8][625] = 16'h0000;
        rom[8][626] = 16'h0000;
        rom[8][627] = 16'h0000;
        rom[8][628] = 16'h0000;
        rom[8][629] = 16'h0000;
        rom[8][630] = 16'h0000;
        rom[8][631] = 16'h0000;
        rom[8][632] = 16'h0000;
        rom[8][633] = 16'h0000;
        rom[8][634] = 16'h0000;
        rom[8][635] = 16'h0000;
        rom[8][636] = 16'h0000;
        rom[8][637] = 16'h0000;
        rom[8][638] = 16'h0000;
        rom[8][639] = 16'h0000;
        rom[8][640] = 16'h0000;
        rom[8][641] = 16'h0000;
        rom[8][642] = 16'h0000;
        rom[8][643] = 16'h0000;
        rom[8][644] = 16'h0000;
        rom[8][645] = 16'h0000;
        rom[8][646] = 16'h0000;
        rom[8][647] = 16'h0000;
        rom[8][648] = 16'h0000;
        rom[8][649] = 16'h0000;
        rom[8][650] = 16'h0000;
        rom[8][651] = 16'h0000;
        rom[8][652] = 16'h0000;
        rom[8][653] = 16'h0000;
        rom[8][654] = 16'h0000;
        rom[8][655] = 16'h0000;
        rom[8][656] = 16'h0000;
        rom[8][657] = 16'h0000;
        rom[8][658] = 16'h0000;
        rom[8][659] = 16'h0000;
        rom[8][660] = 16'h0000;
        rom[8][661] = 16'h0000;
        rom[8][662] = 16'h0000;
        rom[8][663] = 16'h0000;
        rom[8][664] = 16'h0000;
        rom[8][665] = 16'h0000;
        rom[8][666] = 16'h0000;
        rom[8][667] = 16'h0000;
        rom[8][668] = 16'h0000;
        rom[8][669] = 16'h0000;
        rom[8][670] = 16'h0000;
        rom[8][671] = 16'h0000;
        rom[8][672] = 16'h0000;
        rom[8][673] = 16'h0000;
        rom[8][674] = 16'h0000;
        rom[8][675] = 16'h0000;
        rom[8][676] = 16'h0000;
        rom[8][677] = 16'h0000;
        rom[8][678] = 16'h0000;
        rom[8][679] = 16'h0000;
        rom[8][680] = 16'h0000;
        rom[8][681] = 16'h0000;
        rom[8][682] = 16'h0000;
        rom[8][683] = 16'h0000;
        rom[8][684] = 16'h0000;
        rom[8][685] = 16'h0000;
        rom[8][686] = 16'hFEBB;
        rom[8][687] = 16'hFF36;
        rom[8][688] = 16'hFF77;
        rom[8][689] = 16'hFE32;
        rom[8][690] = 16'hFDDB;
        rom[8][691] = 16'hFD9B;
        rom[8][692] = 16'hFE2B;
        rom[8][693] = 16'hFE81;
        rom[8][694] = 16'hFE73;
        rom[8][695] = 16'hFEBB;
        rom[8][696] = 16'hFE1C;
        rom[8][697] = 16'hFDF1;
        rom[8][698] = 16'hFE65;
        rom[8][699] = 16'hFF12;
        rom[8][700] = 16'hFF27;
        rom[8][701] = 16'hFEFC;
        rom[8][702] = 16'hFECA;
        rom[8][703] = 16'hFEDF;
        rom[8][704] = 16'hFF68;
        rom[8][705] = 16'hFE48;
        rom[8][706] = 16'hFE1C;
        rom[8][707] = 16'hFE6C;
        rom[8][708] = 16'hFF0B;
        rom[8][709] = 16'hFF5A;
        rom[8][710] = 16'hFF85;
        rom[8][711] = 16'hFF85;
        rom[8][712] = 16'hFF70;
        rom[8][713] = 16'hFF70;
        rom[8][714] = 16'hFFA2;
        rom[8][715] = 16'hFFC6;
        rom[8][716] = 16'hFF8D;
        rom[8][717] = 16'hFF36;
        rom[8][718] = 16'h0000;
        rom[8][719] = 16'h0000;
        rom[8][720] = 16'h0000;
        rom[8][721] = 16'h0000;
        rom[8][722] = 16'h0000;
        rom[8][723] = 16'h0000;
        rom[8][724] = 16'h0000;
        rom[8][725] = 16'h0000;
        rom[8][726] = 16'h0000;
        rom[8][727] = 16'h0000;
        rom[8][728] = 16'h0000;
        rom[8][729] = 16'h0000;
        rom[8][730] = 16'h0000;
        rom[8][731] = 16'h0000;
        rom[8][732] = 16'h0000;
        rom[8][733] = 16'h0000;
        rom[8][734] = 16'h0000;
        rom[8][735] = 16'h0000;
        rom[8][736] = 16'h0000;
        rom[8][737] = 16'h0000;
        rom[8][738] = 16'h0000;
        rom[8][739] = 16'h0000;
        rom[8][740] = 16'h0000;
        rom[8][741] = 16'h0000;
        rom[8][742] = 16'h0000;
        rom[8][743] = 16'h0000;
        rom[8][744] = 16'h0000;
        rom[8][745] = 16'h0000;
        rom[8][746] = 16'h0000;
        rom[8][747] = 16'h0000;
        rom[8][748] = 16'h0000;
        rom[8][749] = 16'h0000;
        rom[8][750] = 16'h0000;
        rom[8][751] = 16'h0000;
        rom[8][752] = 16'h0000;
        rom[8][753] = 16'h0000;
        rom[8][754] = 16'h0000;
        rom[8][755] = 16'h0000;
        rom[8][756] = 16'h0000;
        rom[8][757] = 16'h0000;
        rom[8][758] = 16'h0000;
        rom[8][759] = 16'h0000;
        rom[8][760] = 16'h0000;
        rom[8][761] = 16'h0000;
        rom[8][762] = 16'h0000;
        rom[8][763] = 16'h0000;
        rom[8][764] = 16'h0000;
        rom[8][765] = 16'h0000;
        rom[8][766] = 16'h0000;
        rom[8][767] = 16'h0000;
        rom[8][768] = 16'h0000;
        rom[8][769] = 16'h0000;
        rom[8][770] = 16'h0000;
        rom[8][771] = 16'h0000;
        rom[8][772] = 16'h0000;
        rom[8][773] = 16'h0000;
        rom[8][774] = 16'h0000;
        rom[8][775] = 16'h0000;
        rom[8][776] = 16'h0000;
        rom[8][777] = 16'h0000;
        rom[8][778] = 16'h0000;
        rom[8][779] = 16'h0000;
        rom[8][780] = 16'h0000;
        rom[8][781] = 16'h0000;
        rom[8][782] = 16'h0000;
        rom[8][783] = 16'h0000;
        rom[8][784] = 16'hFFBF;
        rom[8][785] = 16'h0016;
        rom[8][786] = 16'h003A;
        rom[8][787] = 16'hFF94;
        rom[8][788] = 16'hFF36;
        rom[8][789] = 16'hFF44;
        rom[8][790] = 16'hFF94;
        rom[8][791] = 16'hFF53;
        rom[8][792] = 16'hFF53;
        rom[8][793] = 16'hFFA2;
        rom[8][794] = 16'hFFA2;
        rom[8][795] = 16'hFFB1;
        rom[8][796] = 16'h0016;
        rom[8][797] = 16'h004F;
        rom[8][798] = 16'h001D;
        rom[8][799] = 16'hFFF2;
        rom[8][800] = 16'hFFB8;
        rom[8][801] = 16'hFF85;
        rom[8][802] = 16'hFFA2;
        rom[8][803] = 16'hFF77;
        rom[8][804] = 16'hFF8D;
        rom[8][805] = 16'hFFA9;
        rom[8][806] = 16'h002B;
        rom[8][807] = 16'h0024;
        rom[8][808] = 16'hFFF2;
        rom[8][809] = 16'h0024;
        rom[8][810] = 16'hFFEA;
        rom[8][811] = 16'hFF5A;
        rom[8][812] = 16'hFF77;
        rom[8][813] = 16'hFFA9;
        rom[8][814] = 16'hFF9B;
        rom[8][815] = 16'hFFBF;
        rom[8][816] = 16'h0000;
        rom[8][817] = 16'h0000;
        rom[8][818] = 16'h0000;
        rom[8][819] = 16'h0000;
        rom[8][820] = 16'h0000;
        rom[8][821] = 16'h0000;
        rom[8][822] = 16'h0000;
        rom[8][823] = 16'h0000;
        rom[8][824] = 16'h0000;
        rom[8][825] = 16'h0000;
        rom[8][826] = 16'h0000;
        rom[8][827] = 16'h0000;
        rom[8][828] = 16'h0000;
        rom[8][829] = 16'h0000;
        rom[8][830] = 16'h0000;
        rom[8][831] = 16'h0000;
        rom[8][832] = 16'h0000;
        rom[8][833] = 16'h0000;
        rom[8][834] = 16'h0000;
        rom[8][835] = 16'h0000;
        rom[8][836] = 16'h0000;
        rom[8][837] = 16'h0000;
        rom[8][838] = 16'h0000;
        rom[8][839] = 16'h0000;
        rom[8][840] = 16'h0000;
        rom[8][841] = 16'h0000;
        rom[8][842] = 16'h0000;
        rom[8][843] = 16'h0000;
        rom[8][844] = 16'h0000;
        rom[8][845] = 16'h0000;
        rom[8][846] = 16'h0000;
        rom[8][847] = 16'h0000;
        rom[8][848] = 16'h0000;
        rom[8][849] = 16'h0000;
        rom[8][850] = 16'h0000;
        rom[8][851] = 16'h0000;
        rom[8][852] = 16'h0000;
        rom[8][853] = 16'h0000;
        rom[8][854] = 16'h0000;
        rom[8][855] = 16'h0000;
        rom[8][856] = 16'h0000;
        rom[8][857] = 16'h0000;
        rom[8][858] = 16'h0000;
        rom[8][859] = 16'h0000;
        rom[8][860] = 16'h0000;
        rom[8][861] = 16'h0000;
        rom[8][862] = 16'h0000;
        rom[8][863] = 16'h0000;
        rom[8][864] = 16'h0000;
        rom[8][865] = 16'h0000;
        rom[8][866] = 16'h0000;
        rom[8][867] = 16'h0000;
        rom[8][868] = 16'h0000;
        rom[8][869] = 16'h0000;
        rom[8][870] = 16'h0000;
        rom[8][871] = 16'h0000;
        rom[8][872] = 16'h0000;
        rom[8][873] = 16'h0000;
        rom[8][874] = 16'h0000;
        rom[8][875] = 16'h0000;
        rom[8][876] = 16'h0000;
        rom[8][877] = 16'h0000;
        rom[8][878] = 16'h0000;
        rom[8][879] = 16'h0000;
        rom[8][880] = 16'h0000;
        rom[8][881] = 16'h0000;
        rom[8][882] = 16'h0024;
        rom[8][883] = 16'h0024;
        rom[8][884] = 16'h004F;
        rom[8][885] = 16'h012F;
        rom[8][886] = 16'h0119;
        rom[8][887] = 16'h013E;
        rom[8][888] = 16'h0128;
        rom[8][889] = 16'h00CA;
        rom[8][890] = 16'h0121;
        rom[8][891] = 16'h00E0;
        rom[8][892] = 16'h01C7;
        rom[8][893] = 16'h0208;
        rom[8][894] = 16'h0200;
        rom[8][895] = 16'h0145;
        rom[8][896] = 16'h00EE;
        rom[8][897] = 16'h00EE;
        rom[8][898] = 16'h00E7;
        rom[8][899] = 16'h00B4;
        rom[8][900] = 16'h00D1;
        rom[8][901] = 16'h0112;
        rom[8][902] = 16'h0119;
        rom[8][903] = 16'h010B;
        rom[8][904] = 16'h00FD;
        rom[8][905] = 16'h00E0;
        rom[8][906] = 16'h004F;
        rom[8][907] = 16'h005E;
        rom[8][908] = 16'h003A;
        rom[8][909] = 16'hFFDC;
        rom[8][910] = 16'hFFCD;
        rom[8][911] = 16'h0007;
        rom[8][912] = 16'hFFF9;
        rom[8][913] = 16'h005E;
        rom[8][914] = 16'h0000;
        rom[8][915] = 16'h0000;
        rom[8][916] = 16'h0000;
        rom[8][917] = 16'h0000;
        rom[8][918] = 16'h0000;
        rom[8][919] = 16'h0000;
        rom[8][920] = 16'h0000;
        rom[8][921] = 16'h0000;
        rom[8][922] = 16'h0000;
        rom[8][923] = 16'h0000;
        rom[8][924] = 16'h0000;
        rom[8][925] = 16'h0000;
        rom[8][926] = 16'h0000;
        rom[8][927] = 16'h0000;
        rom[8][928] = 16'h0000;
        rom[8][929] = 16'h0000;
        rom[8][930] = 16'h0000;
        rom[8][931] = 16'h0000;
        rom[8][932] = 16'h0000;
        rom[8][933] = 16'h0000;
        rom[8][934] = 16'h0000;
        rom[8][935] = 16'h0000;
        rom[8][936] = 16'h0000;
        rom[8][937] = 16'h0000;
        rom[8][938] = 16'h0000;
        rom[8][939] = 16'h0000;
        rom[8][940] = 16'h0000;
        rom[8][941] = 16'h0000;
        rom[8][942] = 16'h0000;
        rom[8][943] = 16'h0000;
        rom[8][944] = 16'h0000;
        rom[8][945] = 16'h0000;
        rom[8][946] = 16'h0000;
        rom[8][947] = 16'h0000;
        rom[8][948] = 16'h0000;
        rom[8][949] = 16'h0000;
        rom[8][950] = 16'h0000;
        rom[8][951] = 16'h0000;
        rom[8][952] = 16'h0000;
        rom[8][953] = 16'h0000;
        rom[8][954] = 16'h0000;
        rom[8][955] = 16'h0000;
        rom[8][956] = 16'h0000;
        rom[8][957] = 16'h0000;
        rom[8][958] = 16'h0000;
        rom[8][959] = 16'h0000;
        rom[8][960] = 16'h0000;
        rom[8][961] = 16'h0000;
        rom[8][962] = 16'h0000;
        rom[8][963] = 16'h0000;
        rom[8][964] = 16'h0000;
        rom[8][965] = 16'h0000;
        rom[8][966] = 16'h0000;
        rom[8][967] = 16'h0000;
        rom[8][968] = 16'h0000;
        rom[8][969] = 16'h0000;
        rom[8][970] = 16'h0000;
        rom[8][971] = 16'h0000;
        rom[8][972] = 16'h0000;
        rom[8][973] = 16'h0000;
        rom[8][974] = 16'h0000;
        rom[8][975] = 16'h0000;
        rom[8][976] = 16'h0000;
        rom[8][977] = 16'h0000;
        rom[8][978] = 16'h0000;
        rom[8][979] = 16'h0000;
        rom[8][980] = 16'hFF27;
        rom[8][981] = 16'hFF20;
        rom[8][982] = 16'hFF03;
        rom[8][983] = 16'hFDEA;
        rom[8][984] = 16'hFDA2;
        rom[8][985] = 16'hFE32;
        rom[8][986] = 16'hFE56;
        rom[8][987] = 16'hFEAD;
        rom[8][988] = 16'hFFBF;
        rom[8][989] = 16'hFF27;
        rom[8][990] = 16'hFF7E;
        rom[8][991] = 16'hFFCD;
        rom[8][992] = 16'h0000;
        rom[8][993] = 16'hFFE3;
        rom[8][994] = 16'h000E;
        rom[8][995] = 16'h003A;
        rom[8][996] = 16'h0048;
        rom[8][997] = 16'h007B;
        rom[8][998] = 16'h00D1;
        rom[8][999] = 16'hFF68;
        rom[8][1000] = 16'hFF27;
        rom[8][1001] = 16'hFF36;
        rom[8][1002] = 16'hFF68;
        rom[8][1003] = 16'h003A;
        rom[8][1004] = 16'hFFE3;
        rom[8][1005] = 16'hFFA9;
        rom[8][1006] = 16'hFFA9;
        rom[8][1007] = 16'hFFB1;
        rom[8][1008] = 16'hFFD5;
        rom[8][1009] = 16'hFFEA;
        rom[8][1010] = 16'hFF5A;
        rom[8][1011] = 16'hFF9B;
        rom[8][1012] = 16'h0000;
        rom[8][1013] = 16'h0000;
        rom[8][1014] = 16'h0000;
        rom[8][1015] = 16'h0000;
        rom[8][1016] = 16'h0000;
        rom[8][1017] = 16'h0000;
        rom[8][1018] = 16'h0000;
        rom[8][1019] = 16'h0000;
        rom[8][1020] = 16'h0000;
        rom[8][1021] = 16'h0000;
        rom[8][1022] = 16'h0000;
        rom[8][1023] = 16'h0000;
        rom[8][1024] = 16'h0000;
        rom[8][1025] = 16'h0000;
        rom[8][1026] = 16'h0000;
        rom[8][1027] = 16'h0000;
        rom[8][1028] = 16'h0000;
        rom[8][1029] = 16'h0000;
        rom[8][1030] = 16'h0000;
        rom[8][1031] = 16'h0000;
        rom[8][1032] = 16'h0000;
        rom[8][1033] = 16'h0000;
        rom[8][1034] = 16'h0000;
        rom[8][1035] = 16'h0000;
        rom[8][1036] = 16'h0000;
        rom[8][1037] = 16'h0000;
        rom[8][1038] = 16'h0000;
        rom[8][1039] = 16'h0000;
        rom[8][1040] = 16'h0000;
        rom[8][1041] = 16'h0000;
        rom[8][1042] = 16'h0000;
        rom[8][1043] = 16'h0000;
        rom[8][1044] = 16'h0000;
        rom[8][1045] = 16'h0000;
        rom[8][1046] = 16'h0000;
        rom[8][1047] = 16'h0000;
        rom[8][1048] = 16'h0000;
        rom[8][1049] = 16'h0000;
        rom[8][1050] = 16'h0000;
        rom[8][1051] = 16'h0000;
        rom[8][1052] = 16'h0000;
        rom[8][1053] = 16'h0000;
        rom[8][1054] = 16'h0000;
        rom[8][1055] = 16'h0000;
        rom[8][1056] = 16'h0000;
        rom[8][1057] = 16'h0000;
        rom[8][1058] = 16'h0000;
        rom[8][1059] = 16'h0000;
        rom[8][1060] = 16'h0000;
        rom[8][1061] = 16'h0000;
        rom[8][1062] = 16'h0000;
        rom[8][1063] = 16'h0000;
        rom[8][1064] = 16'h0000;
        rom[8][1065] = 16'h0000;
        rom[8][1066] = 16'h0000;
        rom[8][1067] = 16'h0000;
        rom[8][1068] = 16'h0000;
        rom[8][1069] = 16'h0000;
        rom[8][1070] = 16'h0000;
        rom[8][1071] = 16'h0000;
        rom[8][1072] = 16'h0000;
        rom[8][1073] = 16'h0000;
        rom[8][1074] = 16'h0000;
        rom[8][1075] = 16'h0000;
        rom[8][1076] = 16'h0000;
        rom[8][1077] = 16'h0000;
        rom[8][1078] = 16'hFF68;
        rom[8][1079] = 16'hFF4C;
        rom[8][1080] = 16'hFF3D;
        rom[8][1081] = 16'hFF70;
        rom[8][1082] = 16'h0016;
        rom[8][1083] = 16'h00D9;
        rom[8][1084] = 16'h0104;
        rom[8][1085] = 16'h0104;
        rom[8][1086] = 16'h0136;
        rom[8][1087] = 16'hFFA9;
        rom[8][1088] = 16'hFF4C;
        rom[8][1089] = 16'hFF77;
        rom[8][1090] = 16'hFFC6;
        rom[8][1091] = 16'h0000;
        rom[8][1092] = 16'h0048;
        rom[8][1093] = 16'h00AD;
        rom[8][1094] = 16'h00A6;
        rom[8][1095] = 16'h00B4;
        rom[8][1096] = 16'h0090;
        rom[8][1097] = 16'h003A;
        rom[8][1098] = 16'h0033;
        rom[8][1099] = 16'hFFC6;
        rom[8][1100] = 16'hFF4C;
        rom[8][1101] = 16'hFFBF;
        rom[8][1102] = 16'hFF9B;
        rom[8][1103] = 16'hFF77;
        rom[8][1104] = 16'hFF85;
        rom[8][1105] = 16'hFFD5;
        rom[8][1106] = 16'h0041;
        rom[8][1107] = 16'h000E;
        rom[8][1108] = 16'hFF27;
        rom[8][1109] = 16'hFEE7;
        rom[8][1110] = 16'h0000;
        rom[8][1111] = 16'h0000;
        rom[8][1112] = 16'h0000;
        rom[8][1113] = 16'h0000;
        rom[8][1114] = 16'h0000;
        rom[8][1115] = 16'h0000;
        rom[8][1116] = 16'h0000;
        rom[8][1117] = 16'h0000;
        rom[8][1118] = 16'h0000;
        rom[8][1119] = 16'h0000;
        rom[8][1120] = 16'h0000;
        rom[8][1121] = 16'h0000;
        rom[8][1122] = 16'h0000;
        rom[8][1123] = 16'h0000;
        rom[8][1124] = 16'h0000;
        rom[8][1125] = 16'h0000;
        rom[8][1126] = 16'h0000;
        rom[8][1127] = 16'h0000;
        rom[8][1128] = 16'h0000;
        rom[8][1129] = 16'h0000;
        rom[8][1130] = 16'h0000;
        rom[8][1131] = 16'h0000;
        rom[8][1132] = 16'h0000;
        rom[8][1133] = 16'h0000;
        rom[8][1134] = 16'h0000;
        rom[8][1135] = 16'h0000;
        rom[8][1136] = 16'h0000;
        rom[8][1137] = 16'h0000;
        rom[8][1138] = 16'h0000;
        rom[8][1139] = 16'h0000;
        rom[8][1140] = 16'h0000;
        rom[8][1141] = 16'h0000;
        rom[8][1142] = 16'h0000;
        rom[8][1143] = 16'h0000;
        rom[8][1144] = 16'h0000;
        rom[8][1145] = 16'h0000;
        rom[8][1146] = 16'h0000;
        rom[8][1147] = 16'h0000;
        rom[8][1148] = 16'h0000;
        rom[8][1149] = 16'h0000;
        rom[8][1150] = 16'h0000;
        rom[8][1151] = 16'h0000;
        rom[8][1152] = 16'h0000;
        rom[8][1153] = 16'h0000;
        rom[8][1154] = 16'h0000;
        rom[8][1155] = 16'h0000;
        rom[8][1156] = 16'h0000;
        rom[8][1157] = 16'h0000;
        rom[8][1158] = 16'h0000;
        rom[8][1159] = 16'h0000;
        rom[8][1160] = 16'h0000;
        rom[8][1161] = 16'h0000;
        rom[8][1162] = 16'h0000;
        rom[8][1163] = 16'h0000;
        rom[8][1164] = 16'h0000;
        rom[8][1165] = 16'h0000;
        rom[8][1166] = 16'h0000;
        rom[8][1167] = 16'h0000;
        rom[8][1168] = 16'h0000;
        rom[8][1169] = 16'h0000;
        rom[8][1170] = 16'h0000;
        rom[8][1171] = 16'h0000;
        rom[8][1172] = 16'h0000;
        rom[8][1173] = 16'h0000;
        rom[8][1174] = 16'h0000;
        rom[8][1175] = 16'h0000;
        rom[8][1176] = 16'h0128;
        rom[8][1177] = 16'h00BC;
        rom[8][1178] = 16'h00BC;
        rom[8][1179] = 16'h010B;
        rom[8][1180] = 16'h00EE;
        rom[8][1181] = 16'h0119;
        rom[8][1182] = 16'h010B;
        rom[8][1183] = 16'h00AD;
        rom[8][1184] = 16'h00A6;
        rom[8][1185] = 16'h006C;
        rom[8][1186] = 16'hFFE3;
        rom[8][1187] = 16'hFF94;
        rom[8][1188] = 16'hFF4C;
        rom[8][1189] = 16'hFECA;
        rom[8][1190] = 16'hFEDF;
        rom[8][1191] = 16'hFEF5;
        rom[8][1192] = 16'hFF27;
        rom[8][1193] = 16'hFF8D;
        rom[8][1194] = 16'h002B;
        rom[8][1195] = 16'h0098;
        rom[8][1196] = 16'h0082;
        rom[8][1197] = 16'h0065;
        rom[8][1198] = 16'h0041;
        rom[8][1199] = 16'h0090;
        rom[8][1200] = 16'h004F;
        rom[8][1201] = 16'h0016;
        rom[8][1202] = 16'hFFEA;
        rom[8][1203] = 16'h0065;
        rom[8][1204] = 16'h00E7;
        rom[8][1205] = 16'h00B4;
        rom[8][1206] = 16'h0016;
        rom[8][1207] = 16'hFFC6;
        rom[8][1208] = 16'h0000;
        rom[8][1209] = 16'h0000;
        rom[8][1210] = 16'h0000;
        rom[8][1211] = 16'h0000;
        rom[8][1212] = 16'h0000;
        rom[8][1213] = 16'h0000;
        rom[8][1214] = 16'h0000;
        rom[8][1215] = 16'h0000;
        rom[8][1216] = 16'h0000;
        rom[8][1217] = 16'h0000;
        rom[8][1218] = 16'h0000;
        rom[8][1219] = 16'h0000;
        rom[8][1220] = 16'h0000;
        rom[8][1221] = 16'h0000;
        rom[8][1222] = 16'h0000;
        rom[8][1223] = 16'h0000;
        rom[8][1224] = 16'h0000;
        rom[8][1225] = 16'h0000;
        rom[8][1226] = 16'h0000;
        rom[8][1227] = 16'h0000;
        rom[8][1228] = 16'h0000;
        rom[8][1229] = 16'h0000;
        rom[8][1230] = 16'h0000;
        rom[8][1231] = 16'h0000;
        rom[8][1232] = 16'h0000;
        rom[8][1233] = 16'h0000;
        rom[8][1234] = 16'h0000;
        rom[8][1235] = 16'h0000;
        rom[8][1236] = 16'h0000;
        rom[8][1237] = 16'h0000;
        rom[8][1238] = 16'h0000;
        rom[8][1239] = 16'h0000;
        rom[8][1240] = 16'h0000;
        rom[8][1241] = 16'h0000;
        rom[8][1242] = 16'h0000;
        rom[8][1243] = 16'h0000;
        rom[8][1244] = 16'h0000;
        rom[8][1245] = 16'h0000;
        rom[8][1246] = 16'h0000;
        rom[8][1247] = 16'h0000;
        rom[8][1248] = 16'h0000;
        rom[8][1249] = 16'h0000;
        rom[8][1250] = 16'h0000;
        rom[8][1251] = 16'h0000;
        rom[8][1252] = 16'h0000;
        rom[8][1253] = 16'h0000;
        rom[8][1254] = 16'h0000;
        rom[8][1255] = 16'h0000;
        rom[8][1256] = 16'h0000;
        rom[8][1257] = 16'h0000;
        rom[8][1258] = 16'h0000;
        rom[8][1259] = 16'h0000;
        rom[8][1260] = 16'h0000;
        rom[8][1261] = 16'h0000;
        rom[8][1262] = 16'h0000;
        rom[8][1263] = 16'h0000;
        rom[8][1264] = 16'h0000;
        rom[8][1265] = 16'h0000;
        rom[8][1266] = 16'h0000;
        rom[8][1267] = 16'h0000;
        rom[8][1268] = 16'h0000;
        rom[8][1269] = 16'h0000;
        rom[8][1270] = 16'h0000;
        rom[8][1271] = 16'h0000;
        rom[8][1272] = 16'h0000;
        rom[8][1273] = 16'h0000;
        rom[9][0] = 16'h0073;
        rom[9][1] = 16'h007B;
        rom[9][2] = 16'h006C;
        rom[9][3] = 16'h004F;
        rom[9][4] = 16'h0024;
        rom[9][5] = 16'h000E;
        rom[9][6] = 16'hFFF2;
        rom[9][7] = 16'hFFD5;
        rom[9][8] = 16'hFFB1;
        rom[9][9] = 16'hFF9B;
        rom[9][10] = 16'hFF7E;
        rom[9][11] = 16'hFF61;
        rom[9][12] = 16'hFF53;
        rom[9][13] = 16'hFF4C;
        rom[9][14] = 16'hFFC6;
        rom[9][15] = 16'h0033;
        rom[9][16] = 16'h0073;
        rom[9][17] = 16'h0073;
        rom[9][18] = 16'h006C;
        rom[9][19] = 16'h006C;
        rom[9][20] = 16'h0073;
        rom[9][21] = 16'h0089;
        rom[9][22] = 16'h0098;
        rom[9][23] = 16'h00B4;
        rom[9][24] = 16'h00D1;
        rom[9][25] = 16'h00E7;
        rom[9][26] = 16'h00FD;
        rom[9][27] = 16'h0104;
        rom[9][28] = 16'h0119;
        rom[9][29] = 16'h0112;
        rom[9][30] = 16'h00FD;
        rom[9][31] = 16'h00EE;
        rom[9][32] = 16'h0000;
        rom[9][33] = 16'h0000;
        rom[9][34] = 16'h0000;
        rom[9][35] = 16'h0000;
        rom[9][36] = 16'h0000;
        rom[9][37] = 16'h0000;
        rom[9][38] = 16'h0000;
        rom[9][39] = 16'h0000;
        rom[9][40] = 16'h0000;
        rom[9][41] = 16'h0000;
        rom[9][42] = 16'h0000;
        rom[9][43] = 16'h0000;
        rom[9][44] = 16'h0000;
        rom[9][45] = 16'h0000;
        rom[9][46] = 16'h0000;
        rom[9][47] = 16'h0000;
        rom[9][48] = 16'h0000;
        rom[9][49] = 16'h0000;
        rom[9][50] = 16'h0000;
        rom[9][51] = 16'h0000;
        rom[9][52] = 16'h0000;
        rom[9][53] = 16'h0000;
        rom[9][54] = 16'h0000;
        rom[9][55] = 16'h0000;
        rom[9][56] = 16'h0000;
        rom[9][57] = 16'h0000;
        rom[9][58] = 16'h0000;
        rom[9][59] = 16'h0000;
        rom[9][60] = 16'h0000;
        rom[9][61] = 16'h0000;
        rom[9][62] = 16'h0000;
        rom[9][63] = 16'h0000;
        rom[9][64] = 16'h0000;
        rom[9][65] = 16'h0000;
        rom[9][66] = 16'h0000;
        rom[9][67] = 16'h0000;
        rom[9][68] = 16'h0000;
        rom[9][69] = 16'h0000;
        rom[9][70] = 16'h0000;
        rom[9][71] = 16'h0000;
        rom[9][72] = 16'h0000;
        rom[9][73] = 16'h0000;
        rom[9][74] = 16'h0000;
        rom[9][75] = 16'h0000;
        rom[9][76] = 16'h0000;
        rom[9][77] = 16'h0000;
        rom[9][78] = 16'h0000;
        rom[9][79] = 16'h0000;
        rom[9][80] = 16'h0000;
        rom[9][81] = 16'h0000;
        rom[9][82] = 16'h0000;
        rom[9][83] = 16'h0000;
        rom[9][84] = 16'h0000;
        rom[9][85] = 16'h0000;
        rom[9][86] = 16'h0000;
        rom[9][87] = 16'h0000;
        rom[9][88] = 16'h0000;
        rom[9][89] = 16'h0000;
        rom[9][90] = 16'h0000;
        rom[9][91] = 16'h0000;
        rom[9][92] = 16'h0000;
        rom[9][93] = 16'h0000;
        rom[9][94] = 16'h0000;
        rom[9][95] = 16'h0000;
        rom[9][96] = 16'h0000;
        rom[9][97] = 16'h0000;
        rom[9][98] = 16'h0089;
        rom[9][99] = 16'h006C;
        rom[9][100] = 16'h004F;
        rom[9][101] = 16'h0048;
        rom[9][102] = 16'h0033;
        rom[9][103] = 16'h0024;
        rom[9][104] = 16'h0024;
        rom[9][105] = 16'h000E;
        rom[9][106] = 16'hFFE3;
        rom[9][107] = 16'hFFDC;
        rom[9][108] = 16'hFFCD;
        rom[9][109] = 16'hFFB1;
        rom[9][110] = 16'hFF7E;
        rom[9][111] = 16'hFF53;
        rom[9][112] = 16'h00BC;
        rom[9][113] = 16'h01BF;
        rom[9][114] = 16'h0225;
        rom[9][115] = 16'h023A;
        rom[9][116] = 16'h0225;
        rom[9][117] = 16'h0208;
        rom[9][118] = 16'h01E4;
        rom[9][119] = 16'h01CE;
        rom[9][120] = 16'h01B8;
        rom[9][121] = 16'h01CE;
        rom[9][122] = 16'h01EB;
        rom[9][123] = 16'h01E4;
        rom[9][124] = 16'h01D5;
        rom[9][125] = 16'h01AA;
        rom[9][126] = 16'h018D;
        rom[9][127] = 16'h0177;
        rom[9][128] = 16'h0145;
        rom[9][129] = 16'h012F;
        rom[9][130] = 16'h0000;
        rom[9][131] = 16'h0000;
        rom[9][132] = 16'h0000;
        rom[9][133] = 16'h0000;
        rom[9][134] = 16'h0000;
        rom[9][135] = 16'h0000;
        rom[9][136] = 16'h0000;
        rom[9][137] = 16'h0000;
        rom[9][138] = 16'h0000;
        rom[9][139] = 16'h0000;
        rom[9][140] = 16'h0000;
        rom[9][141] = 16'h0000;
        rom[9][142] = 16'h0000;
        rom[9][143] = 16'h0000;
        rom[9][144] = 16'h0000;
        rom[9][145] = 16'h0000;
        rom[9][146] = 16'h0000;
        rom[9][147] = 16'h0000;
        rom[9][148] = 16'h0000;
        rom[9][149] = 16'h0000;
        rom[9][150] = 16'h0000;
        rom[9][151] = 16'h0000;
        rom[9][152] = 16'h0000;
        rom[9][153] = 16'h0000;
        rom[9][154] = 16'h0000;
        rom[9][155] = 16'h0000;
        rom[9][156] = 16'h0000;
        rom[9][157] = 16'h0000;
        rom[9][158] = 16'h0000;
        rom[9][159] = 16'h0000;
        rom[9][160] = 16'h0000;
        rom[9][161] = 16'h0000;
        rom[9][162] = 16'h0000;
        rom[9][163] = 16'h0000;
        rom[9][164] = 16'h0000;
        rom[9][165] = 16'h0000;
        rom[9][166] = 16'h0000;
        rom[9][167] = 16'h0000;
        rom[9][168] = 16'h0000;
        rom[9][169] = 16'h0000;
        rom[9][170] = 16'h0000;
        rom[9][171] = 16'h0000;
        rom[9][172] = 16'h0000;
        rom[9][173] = 16'h0000;
        rom[9][174] = 16'h0000;
        rom[9][175] = 16'h0000;
        rom[9][176] = 16'h0000;
        rom[9][177] = 16'h0000;
        rom[9][178] = 16'h0000;
        rom[9][179] = 16'h0000;
        rom[9][180] = 16'h0000;
        rom[9][181] = 16'h0000;
        rom[9][182] = 16'h0000;
        rom[9][183] = 16'h0000;
        rom[9][184] = 16'h0000;
        rom[9][185] = 16'h0000;
        rom[9][186] = 16'h0000;
        rom[9][187] = 16'h0000;
        rom[9][188] = 16'h0000;
        rom[9][189] = 16'h0000;
        rom[9][190] = 16'h0000;
        rom[9][191] = 16'h0000;
        rom[9][192] = 16'h0000;
        rom[9][193] = 16'h0000;
        rom[9][194] = 16'h0000;
        rom[9][195] = 16'h0000;
        rom[9][196] = 16'hFE39;
        rom[9][197] = 16'hFE0E;
        rom[9][198] = 16'hFE39;
        rom[9][199] = 16'hFE7A;
        rom[9][200] = 16'hFEA6;
        rom[9][201] = 16'hFEDF;
        rom[9][202] = 16'hFF12;
        rom[9][203] = 16'hFF20;
        rom[9][204] = 16'hFF20;
        rom[9][205] = 16'hFF3D;
        rom[9][206] = 16'hFF7E;
        rom[9][207] = 16'hFFA2;
        rom[9][208] = 16'hFF94;
        rom[9][209] = 16'hFF9B;
        rom[9][210] = 16'h00EE;
        rom[9][211] = 16'h0121;
        rom[9][212] = 16'h0112;
        rom[9][213] = 16'h0136;
        rom[9][214] = 16'h015A;
        rom[9][215] = 16'h014C;
        rom[9][216] = 16'h012F;
        rom[9][217] = 16'h0121;
        rom[9][218] = 16'h0104;
        rom[9][219] = 16'h00E0;
        rom[9][220] = 16'h00E0;
        rom[9][221] = 16'h00D9;
        rom[9][222] = 16'h00E7;
        rom[9][223] = 16'h00BC;
        rom[9][224] = 16'h007B;
        rom[9][225] = 16'h0016;
        rom[9][226] = 16'hFF61;
        rom[9][227] = 16'hFEFC;
        rom[9][228] = 16'h0000;
        rom[9][229] = 16'h0000;
        rom[9][230] = 16'h0000;
        rom[9][231] = 16'h0000;
        rom[9][232] = 16'h0000;
        rom[9][233] = 16'h0000;
        rom[9][234] = 16'h0000;
        rom[9][235] = 16'h0000;
        rom[9][236] = 16'h0000;
        rom[9][237] = 16'h0000;
        rom[9][238] = 16'h0000;
        rom[9][239] = 16'h0000;
        rom[9][240] = 16'h0000;
        rom[9][241] = 16'h0000;
        rom[9][242] = 16'h0000;
        rom[9][243] = 16'h0000;
        rom[9][244] = 16'h0000;
        rom[9][245] = 16'h0000;
        rom[9][246] = 16'h0000;
        rom[9][247] = 16'h0000;
        rom[9][248] = 16'h0000;
        rom[9][249] = 16'h0000;
        rom[9][250] = 16'h0000;
        rom[9][251] = 16'h0000;
        rom[9][252] = 16'h0000;
        rom[9][253] = 16'h0000;
        rom[9][254] = 16'h0000;
        rom[9][255] = 16'h0000;
        rom[9][256] = 16'h0000;
        rom[9][257] = 16'h0000;
        rom[9][258] = 16'h0000;
        rom[9][259] = 16'h0000;
        rom[9][260] = 16'h0000;
        rom[9][261] = 16'h0000;
        rom[9][262] = 16'h0000;
        rom[9][263] = 16'h0000;
        rom[9][264] = 16'h0000;
        rom[9][265] = 16'h0000;
        rom[9][266] = 16'h0000;
        rom[9][267] = 16'h0000;
        rom[9][268] = 16'h0000;
        rom[9][269] = 16'h0000;
        rom[9][270] = 16'h0000;
        rom[9][271] = 16'h0000;
        rom[9][272] = 16'h0000;
        rom[9][273] = 16'h0000;
        rom[9][274] = 16'h0000;
        rom[9][275] = 16'h0000;
        rom[9][276] = 16'h0000;
        rom[9][277] = 16'h0000;
        rom[9][278] = 16'h0000;
        rom[9][279] = 16'h0000;
        rom[9][280] = 16'h0000;
        rom[9][281] = 16'h0000;
        rom[9][282] = 16'h0000;
        rom[9][283] = 16'h0000;
        rom[9][284] = 16'h0000;
        rom[9][285] = 16'h0000;
        rom[9][286] = 16'h0000;
        rom[9][287] = 16'h0000;
        rom[9][288] = 16'h0000;
        rom[9][289] = 16'h0000;
        rom[9][290] = 16'h0000;
        rom[9][291] = 16'h0000;
        rom[9][292] = 16'h0000;
        rom[9][293] = 16'h0000;
        rom[9][294] = 16'hFED8;
        rom[9][295] = 16'hFF5A;
        rom[9][296] = 16'hFFB8;
        rom[9][297] = 16'hFF9B;
        rom[9][298] = 16'hFF5A;
        rom[9][299] = 16'hFF7E;
        rom[9][300] = 16'hFF8D;
        rom[9][301] = 16'hFFA2;
        rom[9][302] = 16'hFF94;
        rom[9][303] = 16'hFF70;
        rom[9][304] = 16'hFFA9;
        rom[9][305] = 16'hFFB8;
        rom[9][306] = 16'hFF7E;
        rom[9][307] = 16'hFF8D;
        rom[9][308] = 16'h0007;
        rom[9][309] = 16'hFFCD;
        rom[9][310] = 16'hFFEA;
        rom[9][311] = 16'hFFDC;
        rom[9][312] = 16'h0024;
        rom[9][313] = 16'h005E;
        rom[9][314] = 16'h00A6;
        rom[9][315] = 16'h00D9;
        rom[9][316] = 16'h00C3;
        rom[9][317] = 16'h0090;
        rom[9][318] = 16'h00A6;
        rom[9][319] = 16'h0128;
        rom[9][320] = 16'h0177;
        rom[9][321] = 16'h0194;
        rom[9][322] = 16'h01C7;
        rom[9][323] = 16'h018D;
        rom[9][324] = 16'h010B;
        rom[9][325] = 16'h00EE;
        rom[9][326] = 16'h0000;
        rom[9][327] = 16'h0000;
        rom[9][328] = 16'h0000;
        rom[9][329] = 16'h0000;
        rom[9][330] = 16'h0000;
        rom[9][331] = 16'h0000;
        rom[9][332] = 16'h0000;
        rom[9][333] = 16'h0000;
        rom[9][334] = 16'h0000;
        rom[9][335] = 16'h0000;
        rom[9][336] = 16'h0000;
        rom[9][337] = 16'h0000;
        rom[9][338] = 16'h0000;
        rom[9][339] = 16'h0000;
        rom[9][340] = 16'h0000;
        rom[9][341] = 16'h0000;
        rom[9][342] = 16'h0000;
        rom[9][343] = 16'h0000;
        rom[9][344] = 16'h0000;
        rom[9][345] = 16'h0000;
        rom[9][346] = 16'h0000;
        rom[9][347] = 16'h0000;
        rom[9][348] = 16'h0000;
        rom[9][349] = 16'h0000;
        rom[9][350] = 16'h0000;
        rom[9][351] = 16'h0000;
        rom[9][352] = 16'h0000;
        rom[9][353] = 16'h0000;
        rom[9][354] = 16'h0000;
        rom[9][355] = 16'h0000;
        rom[9][356] = 16'h0000;
        rom[9][357] = 16'h0000;
        rom[9][358] = 16'h0000;
        rom[9][359] = 16'h0000;
        rom[9][360] = 16'h0000;
        rom[9][361] = 16'h0000;
        rom[9][362] = 16'h0000;
        rom[9][363] = 16'h0000;
        rom[9][364] = 16'h0000;
        rom[9][365] = 16'h0000;
        rom[9][366] = 16'h0000;
        rom[9][367] = 16'h0000;
        rom[9][368] = 16'h0000;
        rom[9][369] = 16'h0000;
        rom[9][370] = 16'h0000;
        rom[9][371] = 16'h0000;
        rom[9][372] = 16'h0000;
        rom[9][373] = 16'h0000;
        rom[9][374] = 16'h0000;
        rom[9][375] = 16'h0000;
        rom[9][376] = 16'h0000;
        rom[9][377] = 16'h0000;
        rom[9][378] = 16'h0000;
        rom[9][379] = 16'h0000;
        rom[9][380] = 16'h0000;
        rom[9][381] = 16'h0000;
        rom[9][382] = 16'h0000;
        rom[9][383] = 16'h0000;
        rom[9][384] = 16'h0000;
        rom[9][385] = 16'h0000;
        rom[9][386] = 16'h0000;
        rom[9][387] = 16'h0000;
        rom[9][388] = 16'h0000;
        rom[9][389] = 16'h0000;
        rom[9][390] = 16'h0000;
        rom[9][391] = 16'h0000;
        rom[9][392] = 16'h0041;
        rom[9][393] = 16'h0082;
        rom[9][394] = 16'h00BC;
        rom[9][395] = 16'h00CA;
        rom[9][396] = 16'h00E7;
        rom[9][397] = 16'h00CA;
        rom[9][398] = 16'h00BC;
        rom[9][399] = 16'h00C3;
        rom[9][400] = 16'h00C3;
        rom[9][401] = 16'h00D9;
        rom[9][402] = 16'h00EE;
        rom[9][403] = 16'h00CA;
        rom[9][404] = 16'h00AD;
        rom[9][405] = 16'h00BC;
        rom[9][406] = 16'h003A;
        rom[9][407] = 16'hFF85;
        rom[9][408] = 16'hFF36;
        rom[9][409] = 16'hFF12;
        rom[9][410] = 16'hFF53;
        rom[9][411] = 16'hFF9B;
        rom[9][412] = 16'hFFEA;
        rom[9][413] = 16'h0024;
        rom[9][414] = 16'h0033;
        rom[9][415] = 16'h001D;
        rom[9][416] = 16'h0041;
        rom[9][417] = 16'h0082;
        rom[9][418] = 16'h0104;
        rom[9][419] = 16'h0169;
        rom[9][420] = 16'h00D1;
        rom[9][421] = 16'h00A6;
        rom[9][422] = 16'h0145;
        rom[9][423] = 16'h0162;
        rom[9][424] = 16'h0000;
        rom[9][425] = 16'h0000;
        rom[9][426] = 16'h0000;
        rom[9][427] = 16'h0000;
        rom[9][428] = 16'h0000;
        rom[9][429] = 16'h0000;
        rom[9][430] = 16'h0000;
        rom[9][431] = 16'h0000;
        rom[9][432] = 16'h0000;
        rom[9][433] = 16'h0000;
        rom[9][434] = 16'h0000;
        rom[9][435] = 16'h0000;
        rom[9][436] = 16'h0000;
        rom[9][437] = 16'h0000;
        rom[9][438] = 16'h0000;
        rom[9][439] = 16'h0000;
        rom[9][440] = 16'h0000;
        rom[9][441] = 16'h0000;
        rom[9][442] = 16'h0000;
        rom[9][443] = 16'h0000;
        rom[9][444] = 16'h0000;
        rom[9][445] = 16'h0000;
        rom[9][446] = 16'h0000;
        rom[9][447] = 16'h0000;
        rom[9][448] = 16'h0000;
        rom[9][449] = 16'h0000;
        rom[9][450] = 16'h0000;
        rom[9][451] = 16'h0000;
        rom[9][452] = 16'h0000;
        rom[9][453] = 16'h0000;
        rom[9][454] = 16'h0000;
        rom[9][455] = 16'h0000;
        rom[9][456] = 16'h0000;
        rom[9][457] = 16'h0000;
        rom[9][458] = 16'h0000;
        rom[9][459] = 16'h0000;
        rom[9][460] = 16'h0000;
        rom[9][461] = 16'h0000;
        rom[9][462] = 16'h0000;
        rom[9][463] = 16'h0000;
        rom[9][464] = 16'h0000;
        rom[9][465] = 16'h0000;
        rom[9][466] = 16'h0000;
        rom[9][467] = 16'h0000;
        rom[9][468] = 16'h0000;
        rom[9][469] = 16'h0000;
        rom[9][470] = 16'h0000;
        rom[9][471] = 16'h0000;
        rom[9][472] = 16'h0000;
        rom[9][473] = 16'h0000;
        rom[9][474] = 16'h0000;
        rom[9][475] = 16'h0000;
        rom[9][476] = 16'h0000;
        rom[9][477] = 16'h0000;
        rom[9][478] = 16'h0000;
        rom[9][479] = 16'h0000;
        rom[9][480] = 16'h0000;
        rom[9][481] = 16'h0000;
        rom[9][482] = 16'h0000;
        rom[9][483] = 16'h0000;
        rom[9][484] = 16'h0000;
        rom[9][485] = 16'h0000;
        rom[9][486] = 16'h0000;
        rom[9][487] = 16'h0000;
        rom[9][488] = 16'h0000;
        rom[9][489] = 16'h0000;
        rom[9][490] = 16'hFFCD;
        rom[9][491] = 16'hFF7E;
        rom[9][492] = 16'hFF8D;
        rom[9][493] = 16'hFFB1;
        rom[9][494] = 16'h0024;
        rom[9][495] = 16'hFFC6;
        rom[9][496] = 16'hFFC6;
        rom[9][497] = 16'hFFCD;
        rom[9][498] = 16'hFFF9;
        rom[9][499] = 16'h001D;
        rom[9][500] = 16'h0000;
        rom[9][501] = 16'hFFCD;
        rom[9][502] = 16'hFFDC;
        rom[9][503] = 16'h0024;
        rom[9][504] = 16'hFEEE;
        rom[9][505] = 16'hFE0E;
        rom[9][506] = 16'hFDD4;
        rom[9][507] = 16'hFDCD;
        rom[9][508] = 16'hFDDB;
        rom[9][509] = 16'hFDF8;
        rom[9][510] = 16'hFDDB;
        rom[9][511] = 16'hFDF8;
        rom[9][512] = 16'hFE65;
        rom[9][513] = 16'hFE4F;
        rom[9][514] = 16'hFE81;
        rom[9][515] = 16'hFF03;
        rom[9][516] = 16'hFF8D;
        rom[9][517] = 16'h0007;
        rom[9][518] = 16'hFFF9;
        rom[9][519] = 16'hFFCD;
        rom[9][520] = 16'hFFF9;
        rom[9][521] = 16'hFFF2;
        rom[9][522] = 16'h0000;
        rom[9][523] = 16'h0000;
        rom[9][524] = 16'h0000;
        rom[9][525] = 16'h0000;
        rom[9][526] = 16'h0000;
        rom[9][527] = 16'h0000;
        rom[9][528] = 16'h0000;
        rom[9][529] = 16'h0000;
        rom[9][530] = 16'h0000;
        rom[9][531] = 16'h0000;
        rom[9][532] = 16'h0000;
        rom[9][533] = 16'h0000;
        rom[9][534] = 16'h0000;
        rom[9][535] = 16'h0000;
        rom[9][536] = 16'h0000;
        rom[9][537] = 16'h0000;
        rom[9][538] = 16'h0000;
        rom[9][539] = 16'h0000;
        rom[9][540] = 16'h0000;
        rom[9][541] = 16'h0000;
        rom[9][542] = 16'h0000;
        rom[9][543] = 16'h0000;
        rom[9][544] = 16'h0000;
        rom[9][545] = 16'h0000;
        rom[9][546] = 16'h0000;
        rom[9][547] = 16'h0000;
        rom[9][548] = 16'h0000;
        rom[9][549] = 16'h0000;
        rom[9][550] = 16'h0000;
        rom[9][551] = 16'h0000;
        rom[9][552] = 16'h0000;
        rom[9][553] = 16'h0000;
        rom[9][554] = 16'h0000;
        rom[9][555] = 16'h0000;
        rom[9][556] = 16'h0000;
        rom[9][557] = 16'h0000;
        rom[9][558] = 16'h0000;
        rom[9][559] = 16'h0000;
        rom[9][560] = 16'h0000;
        rom[9][561] = 16'h0000;
        rom[9][562] = 16'h0000;
        rom[9][563] = 16'h0000;
        rom[9][564] = 16'h0000;
        rom[9][565] = 16'h0000;
        rom[9][566] = 16'h0000;
        rom[9][567] = 16'h0000;
        rom[9][568] = 16'h0000;
        rom[9][569] = 16'h0000;
        rom[9][570] = 16'h0000;
        rom[9][571] = 16'h0000;
        rom[9][572] = 16'h0000;
        rom[9][573] = 16'h0000;
        rom[9][574] = 16'h0000;
        rom[9][575] = 16'h0000;
        rom[9][576] = 16'h0000;
        rom[9][577] = 16'h0000;
        rom[9][578] = 16'h0000;
        rom[9][579] = 16'h0000;
        rom[9][580] = 16'h0000;
        rom[9][581] = 16'h0000;
        rom[9][582] = 16'h0000;
        rom[9][583] = 16'h0000;
        rom[9][584] = 16'h0000;
        rom[9][585] = 16'h0000;
        rom[9][586] = 16'h0000;
        rom[9][587] = 16'h0000;
        rom[9][588] = 16'h007B;
        rom[9][589] = 16'h006C;
        rom[9][590] = 16'h0082;
        rom[9][591] = 16'h0065;
        rom[9][592] = 16'h005E;
        rom[9][593] = 16'h003A;
        rom[9][594] = 16'h0065;
        rom[9][595] = 16'h00B4;
        rom[9][596] = 16'h00E0;
        rom[9][597] = 16'h00D9;
        rom[9][598] = 16'h00C3;
        rom[9][599] = 16'h0073;
        rom[9][600] = 16'h002B;
        rom[9][601] = 16'h0057;
        rom[9][602] = 16'hFF85;
        rom[9][603] = 16'hFF8D;
        rom[9][604] = 16'hFFB8;
        rom[9][605] = 16'hFFCD;
        rom[9][606] = 16'hFFA9;
        rom[9][607] = 16'hFF61;
        rom[9][608] = 16'hFEFC;
        rom[9][609] = 16'hFEFC;
        rom[9][610] = 16'hFF36;
        rom[9][611] = 16'hFF5A;
        rom[9][612] = 16'hFF9B;
        rom[9][613] = 16'hFFDC;
        rom[9][614] = 16'hFFC6;
        rom[9][615] = 16'hFFE3;
        rom[9][616] = 16'h004F;
        rom[9][617] = 16'h006C;
        rom[9][618] = 16'h002B;
        rom[9][619] = 16'hFFF2;
        rom[9][620] = 16'h0000;
        rom[9][621] = 16'h0000;
        rom[9][622] = 16'h0000;
        rom[9][623] = 16'h0000;
        rom[9][624] = 16'h0000;
        rom[9][625] = 16'h0000;
        rom[9][626] = 16'h0000;
        rom[9][627] = 16'h0000;
        rom[9][628] = 16'h0000;
        rom[9][629] = 16'h0000;
        rom[9][630] = 16'h0000;
        rom[9][631] = 16'h0000;
        rom[9][632] = 16'h0000;
        rom[9][633] = 16'h0000;
        rom[9][634] = 16'h0000;
        rom[9][635] = 16'h0000;
        rom[9][636] = 16'h0000;
        rom[9][637] = 16'h0000;
        rom[9][638] = 16'h0000;
        rom[9][639] = 16'h0000;
        rom[9][640] = 16'h0000;
        rom[9][641] = 16'h0000;
        rom[9][642] = 16'h0000;
        rom[9][643] = 16'h0000;
        rom[9][644] = 16'h0000;
        rom[9][645] = 16'h0000;
        rom[9][646] = 16'h0000;
        rom[9][647] = 16'h0000;
        rom[9][648] = 16'h0000;
        rom[9][649] = 16'h0000;
        rom[9][650] = 16'h0000;
        rom[9][651] = 16'h0000;
        rom[9][652] = 16'h0000;
        rom[9][653] = 16'h0000;
        rom[9][654] = 16'h0000;
        rom[9][655] = 16'h0000;
        rom[9][656] = 16'h0000;
        rom[9][657] = 16'h0000;
        rom[9][658] = 16'h0000;
        rom[9][659] = 16'h0000;
        rom[9][660] = 16'h0000;
        rom[9][661] = 16'h0000;
        rom[9][662] = 16'h0000;
        rom[9][663] = 16'h0000;
        rom[9][664] = 16'h0000;
        rom[9][665] = 16'h0000;
        rom[9][666] = 16'h0000;
        rom[9][667] = 16'h0000;
        rom[9][668] = 16'h0000;
        rom[9][669] = 16'h0000;
        rom[9][670] = 16'h0000;
        rom[9][671] = 16'h0000;
        rom[9][672] = 16'h0000;
        rom[9][673] = 16'h0000;
        rom[9][674] = 16'h0000;
        rom[9][675] = 16'h0000;
        rom[9][676] = 16'h0000;
        rom[9][677] = 16'h0000;
        rom[9][678] = 16'h0000;
        rom[9][679] = 16'h0000;
        rom[9][680] = 16'h0000;
        rom[9][681] = 16'h0000;
        rom[9][682] = 16'h0000;
        rom[9][683] = 16'h0000;
        rom[9][684] = 16'h0000;
        rom[9][685] = 16'h0000;
        rom[9][686] = 16'h0098;
        rom[9][687] = 16'h0041;
        rom[9][688] = 16'h0041;
        rom[9][689] = 16'h0089;
        rom[9][690] = 16'h0090;
        rom[9][691] = 16'h00E0;
        rom[9][692] = 16'h0136;
        rom[9][693] = 16'h0121;
        rom[9][694] = 16'h00FD;
        rom[9][695] = 16'h00BC;
        rom[9][696] = 16'h00AD;
        rom[9][697] = 16'h00D9;
        rom[9][698] = 16'h00F5;
        rom[9][699] = 16'h015A;
        rom[9][700] = 16'h0112;
        rom[9][701] = 16'h0128;
        rom[9][702] = 16'h0104;
        rom[9][703] = 16'h00B4;
        rom[9][704] = 16'h00AD;
        rom[9][705] = 16'h006C;
        rom[9][706] = 16'h0024;
        rom[9][707] = 16'h004F;
        rom[9][708] = 16'h0041;
        rom[9][709] = 16'h002B;
        rom[9][710] = 16'h003A;
        rom[9][711] = 16'hFFCD;
        rom[9][712] = 16'hFF85;
        rom[9][713] = 16'hFF53;
        rom[9][714] = 16'hFF27;
        rom[9][715] = 16'hFEFC;
        rom[9][716] = 16'hFF94;
        rom[9][717] = 16'h0016;
        rom[9][718] = 16'h0000;
        rom[9][719] = 16'h0000;
        rom[9][720] = 16'h0000;
        rom[9][721] = 16'h0000;
        rom[9][722] = 16'h0000;
        rom[9][723] = 16'h0000;
        rom[9][724] = 16'h0000;
        rom[9][725] = 16'h0000;
        rom[9][726] = 16'h0000;
        rom[9][727] = 16'h0000;
        rom[9][728] = 16'h0000;
        rom[9][729] = 16'h0000;
        rom[9][730] = 16'h0000;
        rom[9][731] = 16'h0000;
        rom[9][732] = 16'h0000;
        rom[9][733] = 16'h0000;
        rom[9][734] = 16'h0000;
        rom[9][735] = 16'h0000;
        rom[9][736] = 16'h0000;
        rom[9][737] = 16'h0000;
        rom[9][738] = 16'h0000;
        rom[9][739] = 16'h0000;
        rom[9][740] = 16'h0000;
        rom[9][741] = 16'h0000;
        rom[9][742] = 16'h0000;
        rom[9][743] = 16'h0000;
        rom[9][744] = 16'h0000;
        rom[9][745] = 16'h0000;
        rom[9][746] = 16'h0000;
        rom[9][747] = 16'h0000;
        rom[9][748] = 16'h0000;
        rom[9][749] = 16'h0000;
        rom[9][750] = 16'h0000;
        rom[9][751] = 16'h0000;
        rom[9][752] = 16'h0000;
        rom[9][753] = 16'h0000;
        rom[9][754] = 16'h0000;
        rom[9][755] = 16'h0000;
        rom[9][756] = 16'h0000;
        rom[9][757] = 16'h0000;
        rom[9][758] = 16'h0000;
        rom[9][759] = 16'h0000;
        rom[9][760] = 16'h0000;
        rom[9][761] = 16'h0000;
        rom[9][762] = 16'h0000;
        rom[9][763] = 16'h0000;
        rom[9][764] = 16'h0000;
        rom[9][765] = 16'h0000;
        rom[9][766] = 16'h0000;
        rom[9][767] = 16'h0000;
        rom[9][768] = 16'h0000;
        rom[9][769] = 16'h0000;
        rom[9][770] = 16'h0000;
        rom[9][771] = 16'h0000;
        rom[9][772] = 16'h0000;
        rom[9][773] = 16'h0000;
        rom[9][774] = 16'h0000;
        rom[9][775] = 16'h0000;
        rom[9][776] = 16'h0000;
        rom[9][777] = 16'h0000;
        rom[9][778] = 16'h0000;
        rom[9][779] = 16'h0000;
        rom[9][780] = 16'h0000;
        rom[9][781] = 16'h0000;
        rom[9][782] = 16'h0000;
        rom[9][783] = 16'h0000;
        rom[9][784] = 16'hFFCD;
        rom[9][785] = 16'hFF53;
        rom[9][786] = 16'hFF61;
        rom[9][787] = 16'hFF85;
        rom[9][788] = 16'hFFB8;
        rom[9][789] = 16'h001D;
        rom[9][790] = 16'h002B;
        rom[9][791] = 16'h000E;
        rom[9][792] = 16'hFFEA;
        rom[9][793] = 16'hFFBF;
        rom[9][794] = 16'hFFEA;
        rom[9][795] = 16'h001D;
        rom[9][796] = 16'hFFC6;
        rom[9][797] = 16'hFF85;
        rom[9][798] = 16'hFFB8;
        rom[9][799] = 16'h006C;
        rom[9][800] = 16'h0082;
        rom[9][801] = 16'h003A;
        rom[9][802] = 16'h001D;
        rom[9][803] = 16'h007B;
        rom[9][804] = 16'h0016;
        rom[9][805] = 16'hFFF9;
        rom[9][806] = 16'h0090;
        rom[9][807] = 16'h0065;
        rom[9][808] = 16'h003A;
        rom[9][809] = 16'hFF4C;
        rom[9][810] = 16'hFE32;
        rom[9][811] = 16'hFE15;
        rom[9][812] = 16'hFF12;
        rom[9][813] = 16'hFF61;
        rom[9][814] = 16'hFF77;
        rom[9][815] = 16'h003A;
        rom[9][816] = 16'h0000;
        rom[9][817] = 16'h0000;
        rom[9][818] = 16'h0000;
        rom[9][819] = 16'h0000;
        rom[9][820] = 16'h0000;
        rom[9][821] = 16'h0000;
        rom[9][822] = 16'h0000;
        rom[9][823] = 16'h0000;
        rom[9][824] = 16'h0000;
        rom[9][825] = 16'h0000;
        rom[9][826] = 16'h0000;
        rom[9][827] = 16'h0000;
        rom[9][828] = 16'h0000;
        rom[9][829] = 16'h0000;
        rom[9][830] = 16'h0000;
        rom[9][831] = 16'h0000;
        rom[9][832] = 16'h0000;
        rom[9][833] = 16'h0000;
        rom[9][834] = 16'h0000;
        rom[9][835] = 16'h0000;
        rom[9][836] = 16'h0000;
        rom[9][837] = 16'h0000;
        rom[9][838] = 16'h0000;
        rom[9][839] = 16'h0000;
        rom[9][840] = 16'h0000;
        rom[9][841] = 16'h0000;
        rom[9][842] = 16'h0000;
        rom[9][843] = 16'h0000;
        rom[9][844] = 16'h0000;
        rom[9][845] = 16'h0000;
        rom[9][846] = 16'h0000;
        rom[9][847] = 16'h0000;
        rom[9][848] = 16'h0000;
        rom[9][849] = 16'h0000;
        rom[9][850] = 16'h0000;
        rom[9][851] = 16'h0000;
        rom[9][852] = 16'h0000;
        rom[9][853] = 16'h0000;
        rom[9][854] = 16'h0000;
        rom[9][855] = 16'h0000;
        rom[9][856] = 16'h0000;
        rom[9][857] = 16'h0000;
        rom[9][858] = 16'h0000;
        rom[9][859] = 16'h0000;
        rom[9][860] = 16'h0000;
        rom[9][861] = 16'h0000;
        rom[9][862] = 16'h0000;
        rom[9][863] = 16'h0000;
        rom[9][864] = 16'h0000;
        rom[9][865] = 16'h0000;
        rom[9][866] = 16'h0000;
        rom[9][867] = 16'h0000;
        rom[9][868] = 16'h0000;
        rom[9][869] = 16'h0000;
        rom[9][870] = 16'h0000;
        rom[9][871] = 16'h0000;
        rom[9][872] = 16'h0000;
        rom[9][873] = 16'h0000;
        rom[9][874] = 16'h0000;
        rom[9][875] = 16'h0000;
        rom[9][876] = 16'h0000;
        rom[9][877] = 16'h0000;
        rom[9][878] = 16'h0000;
        rom[9][879] = 16'h0000;
        rom[9][880] = 16'h0000;
        rom[9][881] = 16'h0000;
        rom[9][882] = 16'hFFC6;
        rom[9][883] = 16'hFFB8;
        rom[9][884] = 16'hFFBF;
        rom[9][885] = 16'hFF7E;
        rom[9][886] = 16'hFF36;
        rom[9][887] = 16'hFFD5;
        rom[9][888] = 16'h001D;
        rom[9][889] = 16'h0000;
        rom[9][890] = 16'hFF77;
        rom[9][891] = 16'hFF36;
        rom[9][892] = 16'hFF53;
        rom[9][893] = 16'hFFC6;
        rom[9][894] = 16'h0057;
        rom[9][895] = 16'h007B;
        rom[9][896] = 16'h0024;
        rom[9][897] = 16'hFFE3;
        rom[9][898] = 16'hFF77;
        rom[9][899] = 16'hFF7E;
        rom[9][900] = 16'hFFF2;
        rom[9][901] = 16'h0041;
        rom[9][902] = 16'hFFF2;
        rom[9][903] = 16'h001D;
        rom[9][904] = 16'h0098;
        rom[9][905] = 16'h007B;
        rom[9][906] = 16'h0048;
        rom[9][907] = 16'h002B;
        rom[9][908] = 16'hFF5A;
        rom[9][909] = 16'hFF2F;
        rom[9][910] = 16'hFFD5;
        rom[9][911] = 16'hFFC6;
        rom[9][912] = 16'hFFDC;
        rom[9][913] = 16'h0048;
        rom[9][914] = 16'h0000;
        rom[9][915] = 16'h0000;
        rom[9][916] = 16'h0000;
        rom[9][917] = 16'h0000;
        rom[9][918] = 16'h0000;
        rom[9][919] = 16'h0000;
        rom[9][920] = 16'h0000;
        rom[9][921] = 16'h0000;
        rom[9][922] = 16'h0000;
        rom[9][923] = 16'h0000;
        rom[9][924] = 16'h0000;
        rom[9][925] = 16'h0000;
        rom[9][926] = 16'h0000;
        rom[9][927] = 16'h0000;
        rom[9][928] = 16'h0000;
        rom[9][929] = 16'h0000;
        rom[9][930] = 16'h0000;
        rom[9][931] = 16'h0000;
        rom[9][932] = 16'h0000;
        rom[9][933] = 16'h0000;
        rom[9][934] = 16'h0000;
        rom[9][935] = 16'h0000;
        rom[9][936] = 16'h0000;
        rom[9][937] = 16'h0000;
        rom[9][938] = 16'h0000;
        rom[9][939] = 16'h0000;
        rom[9][940] = 16'h0000;
        rom[9][941] = 16'h0000;
        rom[9][942] = 16'h0000;
        rom[9][943] = 16'h0000;
        rom[9][944] = 16'h0000;
        rom[9][945] = 16'h0000;
        rom[9][946] = 16'h0000;
        rom[9][947] = 16'h0000;
        rom[9][948] = 16'h0000;
        rom[9][949] = 16'h0000;
        rom[9][950] = 16'h0000;
        rom[9][951] = 16'h0000;
        rom[9][952] = 16'h0000;
        rom[9][953] = 16'h0000;
        rom[9][954] = 16'h0000;
        rom[9][955] = 16'h0000;
        rom[9][956] = 16'h0000;
        rom[9][957] = 16'h0000;
        rom[9][958] = 16'h0000;
        rom[9][959] = 16'h0000;
        rom[9][960] = 16'h0000;
        rom[9][961] = 16'h0000;
        rom[9][962] = 16'h0000;
        rom[9][963] = 16'h0000;
        rom[9][964] = 16'h0000;
        rom[9][965] = 16'h0000;
        rom[9][966] = 16'h0000;
        rom[9][967] = 16'h0000;
        rom[9][968] = 16'h0000;
        rom[9][969] = 16'h0000;
        rom[9][970] = 16'h0000;
        rom[9][971] = 16'h0000;
        rom[9][972] = 16'h0000;
        rom[9][973] = 16'h0000;
        rom[9][974] = 16'h0000;
        rom[9][975] = 16'h0000;
        rom[9][976] = 16'h0000;
        rom[9][977] = 16'h0000;
        rom[9][978] = 16'h0000;
        rom[9][979] = 16'h0000;
        rom[9][980] = 16'h0073;
        rom[9][981] = 16'h002B;
        rom[9][982] = 16'hFFBF;
        rom[9][983] = 16'hFFD5;
        rom[9][984] = 16'h0016;
        rom[9][985] = 16'h0033;
        rom[9][986] = 16'h0089;
        rom[9][987] = 16'h004F;
        rom[9][988] = 16'hFFF2;
        rom[9][989] = 16'hFFD5;
        rom[9][990] = 16'hFFB1;
        rom[9][991] = 16'hFFE3;
        rom[9][992] = 16'h0048;
        rom[9][993] = 16'h0065;
        rom[9][994] = 16'hFF7E;
        rom[9][995] = 16'hFF27;
        rom[9][996] = 16'hFEFC;
        rom[9][997] = 16'hFF44;
        rom[9][998] = 16'hFF9B;
        rom[9][999] = 16'hFF85;
        rom[9][1000] = 16'hFF8D;
        rom[9][1001] = 16'hFF7E;
        rom[9][1002] = 16'hFF61;
        rom[9][1003] = 16'hFF77;
        rom[9][1004] = 16'hFFCD;
        rom[9][1005] = 16'h0000;
        rom[9][1006] = 16'h000E;
        rom[9][1007] = 16'hFFCD;
        rom[9][1008] = 16'hFFC6;
        rom[9][1009] = 16'hFFEA;
        rom[9][1010] = 16'hFFD5;
        rom[9][1011] = 16'hFFF9;
        rom[9][1012] = 16'h0000;
        rom[9][1013] = 16'h0000;
        rom[9][1014] = 16'h0000;
        rom[9][1015] = 16'h0000;
        rom[9][1016] = 16'h0000;
        rom[9][1017] = 16'h0000;
        rom[9][1018] = 16'h0000;
        rom[9][1019] = 16'h0000;
        rom[9][1020] = 16'h0000;
        rom[9][1021] = 16'h0000;
        rom[9][1022] = 16'h0000;
        rom[9][1023] = 16'h0000;
        rom[9][1024] = 16'h0000;
        rom[9][1025] = 16'h0000;
        rom[9][1026] = 16'h0000;
        rom[9][1027] = 16'h0000;
        rom[9][1028] = 16'h0000;
        rom[9][1029] = 16'h0000;
        rom[9][1030] = 16'h0000;
        rom[9][1031] = 16'h0000;
        rom[9][1032] = 16'h0000;
        rom[9][1033] = 16'h0000;
        rom[9][1034] = 16'h0000;
        rom[9][1035] = 16'h0000;
        rom[9][1036] = 16'h0000;
        rom[9][1037] = 16'h0000;
        rom[9][1038] = 16'h0000;
        rom[9][1039] = 16'h0000;
        rom[9][1040] = 16'h0000;
        rom[9][1041] = 16'h0000;
        rom[9][1042] = 16'h0000;
        rom[9][1043] = 16'h0000;
        rom[9][1044] = 16'h0000;
        rom[9][1045] = 16'h0000;
        rom[9][1046] = 16'h0000;
        rom[9][1047] = 16'h0000;
        rom[9][1048] = 16'h0000;
        rom[9][1049] = 16'h0000;
        rom[9][1050] = 16'h0000;
        rom[9][1051] = 16'h0000;
        rom[9][1052] = 16'h0000;
        rom[9][1053] = 16'h0000;
        rom[9][1054] = 16'h0000;
        rom[9][1055] = 16'h0000;
        rom[9][1056] = 16'h0000;
        rom[9][1057] = 16'h0000;
        rom[9][1058] = 16'h0000;
        rom[9][1059] = 16'h0000;
        rom[9][1060] = 16'h0000;
        rom[9][1061] = 16'h0000;
        rom[9][1062] = 16'h0000;
        rom[9][1063] = 16'h0000;
        rom[9][1064] = 16'h0000;
        rom[9][1065] = 16'h0000;
        rom[9][1066] = 16'h0000;
        rom[9][1067] = 16'h0000;
        rom[9][1068] = 16'h0000;
        rom[9][1069] = 16'h0000;
        rom[9][1070] = 16'h0000;
        rom[9][1071] = 16'h0000;
        rom[9][1072] = 16'h0000;
        rom[9][1073] = 16'h0000;
        rom[9][1074] = 16'h0000;
        rom[9][1075] = 16'h0000;
        rom[9][1076] = 16'h0000;
        rom[9][1077] = 16'h0000;
        rom[9][1078] = 16'hFFB1;
        rom[9][1079] = 16'hFF27;
        rom[9][1080] = 16'hFEF5;
        rom[9][1081] = 16'hFFCD;
        rom[9][1082] = 16'h002B;
        rom[9][1083] = 16'h0057;
        rom[9][1084] = 16'h0048;
        rom[9][1085] = 16'hFFB1;
        rom[9][1086] = 16'hFF9B;
        rom[9][1087] = 16'hFFA2;
        rom[9][1088] = 16'hFFF9;
        rom[9][1089] = 16'hFFF9;
        rom[9][1090] = 16'h0007;
        rom[9][1091] = 16'hFFE3;
        rom[9][1092] = 16'hFF4C;
        rom[9][1093] = 16'hFF4C;
        rom[9][1094] = 16'hFF12;
        rom[9][1095] = 16'hFEE7;
        rom[9][1096] = 16'hFEB4;
        rom[9][1097] = 16'hFECA;
        rom[9][1098] = 16'hFF5A;
        rom[9][1099] = 16'hFF03;
        rom[9][1100] = 16'hFED1;
        rom[9][1101] = 16'hFF3D;
        rom[9][1102] = 16'hFF8D;
        rom[9][1103] = 16'hFFE3;
        rom[9][1104] = 16'h000E;
        rom[9][1105] = 16'hFFD5;
        rom[9][1106] = 16'h0082;
        rom[9][1107] = 16'h0104;
        rom[9][1108] = 16'h00B4;
        rom[9][1109] = 16'h0121;
        rom[9][1110] = 16'h0000;
        rom[9][1111] = 16'h0000;
        rom[9][1112] = 16'h0000;
        rom[9][1113] = 16'h0000;
        rom[9][1114] = 16'h0000;
        rom[9][1115] = 16'h0000;
        rom[9][1116] = 16'h0000;
        rom[9][1117] = 16'h0000;
        rom[9][1118] = 16'h0000;
        rom[9][1119] = 16'h0000;
        rom[9][1120] = 16'h0000;
        rom[9][1121] = 16'h0000;
        rom[9][1122] = 16'h0000;
        rom[9][1123] = 16'h0000;
        rom[9][1124] = 16'h0000;
        rom[9][1125] = 16'h0000;
        rom[9][1126] = 16'h0000;
        rom[9][1127] = 16'h0000;
        rom[9][1128] = 16'h0000;
        rom[9][1129] = 16'h0000;
        rom[9][1130] = 16'h0000;
        rom[9][1131] = 16'h0000;
        rom[9][1132] = 16'h0000;
        rom[9][1133] = 16'h0000;
        rom[9][1134] = 16'h0000;
        rom[9][1135] = 16'h0000;
        rom[9][1136] = 16'h0000;
        rom[9][1137] = 16'h0000;
        rom[9][1138] = 16'h0000;
        rom[9][1139] = 16'h0000;
        rom[9][1140] = 16'h0000;
        rom[9][1141] = 16'h0000;
        rom[9][1142] = 16'h0000;
        rom[9][1143] = 16'h0000;
        rom[9][1144] = 16'h0000;
        rom[9][1145] = 16'h0000;
        rom[9][1146] = 16'h0000;
        rom[9][1147] = 16'h0000;
        rom[9][1148] = 16'h0000;
        rom[9][1149] = 16'h0000;
        rom[9][1150] = 16'h0000;
        rom[9][1151] = 16'h0000;
        rom[9][1152] = 16'h0000;
        rom[9][1153] = 16'h0000;
        rom[9][1154] = 16'h0000;
        rom[9][1155] = 16'h0000;
        rom[9][1156] = 16'h0000;
        rom[9][1157] = 16'h0000;
        rom[9][1158] = 16'h0000;
        rom[9][1159] = 16'h0000;
        rom[9][1160] = 16'h0000;
        rom[9][1161] = 16'h0000;
        rom[9][1162] = 16'h0000;
        rom[9][1163] = 16'h0000;
        rom[9][1164] = 16'h0000;
        rom[9][1165] = 16'h0000;
        rom[9][1166] = 16'h0000;
        rom[9][1167] = 16'h0000;
        rom[9][1168] = 16'h0000;
        rom[9][1169] = 16'h0000;
        rom[9][1170] = 16'h0000;
        rom[9][1171] = 16'h0000;
        rom[9][1172] = 16'h0000;
        rom[9][1173] = 16'h0000;
        rom[9][1174] = 16'h0000;
        rom[9][1175] = 16'h0000;
        rom[9][1176] = 16'h0000;
        rom[9][1177] = 16'h009F;
        rom[9][1178] = 16'h0098;
        rom[9][1179] = 16'h0057;
        rom[9][1180] = 16'h0057;
        rom[9][1181] = 16'h00D9;
        rom[9][1182] = 16'h00EE;
        rom[9][1183] = 16'h006C;
        rom[9][1184] = 16'h0082;
        rom[9][1185] = 16'h0000;
        rom[9][1186] = 16'hFFB8;
        rom[9][1187] = 16'h000E;
        rom[9][1188] = 16'hFFC6;
        rom[9][1189] = 16'hFFCD;
        rom[9][1190] = 16'hFF53;
        rom[9][1191] = 16'hFF61;
        rom[9][1192] = 16'hFF44;
        rom[9][1193] = 16'hFF44;
        rom[9][1194] = 16'hFF7E;
        rom[9][1195] = 16'hFFA2;
        rom[9][1196] = 16'hFFDC;
        rom[9][1197] = 16'hFFBF;
        rom[9][1198] = 16'hFFBF;
        rom[9][1199] = 16'hFFEA;
        rom[9][1200] = 16'h0089;
        rom[9][1201] = 16'h0119;
        rom[9][1202] = 16'h00C3;
        rom[9][1203] = 16'h0048;
        rom[9][1204] = 16'h005E;
        rom[9][1205] = 16'h00AD;
        rom[9][1206] = 16'h0104;
        rom[9][1207] = 16'h0162;
        rom[9][1208] = 16'h0000;
        rom[9][1209] = 16'h0000;
        rom[9][1210] = 16'h0000;
        rom[9][1211] = 16'h0000;
        rom[9][1212] = 16'h0000;
        rom[9][1213] = 16'h0000;
        rom[9][1214] = 16'h0000;
        rom[9][1215] = 16'h0000;
        rom[9][1216] = 16'h0000;
        rom[9][1217] = 16'h0000;
        rom[9][1218] = 16'h0000;
        rom[9][1219] = 16'h0000;
        rom[9][1220] = 16'h0000;
        rom[9][1221] = 16'h0000;
        rom[9][1222] = 16'h0000;
        rom[9][1223] = 16'h0000;
        rom[9][1224] = 16'h0000;
        rom[9][1225] = 16'h0000;
        rom[9][1226] = 16'h0000;
        rom[9][1227] = 16'h0000;
        rom[9][1228] = 16'h0000;
        rom[9][1229] = 16'h0000;
        rom[9][1230] = 16'h0000;
        rom[9][1231] = 16'h0000;
        rom[9][1232] = 16'h0000;
        rom[9][1233] = 16'h0000;
        rom[9][1234] = 16'h0000;
        rom[9][1235] = 16'h0000;
        rom[9][1236] = 16'h0000;
        rom[9][1237] = 16'h0000;
        rom[9][1238] = 16'h0000;
        rom[9][1239] = 16'h0000;
        rom[9][1240] = 16'h0000;
        rom[9][1241] = 16'h0000;
        rom[9][1242] = 16'h0000;
        rom[9][1243] = 16'h0000;
        rom[9][1244] = 16'h0000;
        rom[9][1245] = 16'h0000;
        rom[9][1246] = 16'h0000;
        rom[9][1247] = 16'h0000;
        rom[9][1248] = 16'h0000;
        rom[9][1249] = 16'h0000;
        rom[9][1250] = 16'h0000;
        rom[9][1251] = 16'h0000;
        rom[9][1252] = 16'h0000;
        rom[9][1253] = 16'h0000;
        rom[9][1254] = 16'h0000;
        rom[9][1255] = 16'h0000;
        rom[9][1256] = 16'h0000;
        rom[9][1257] = 16'h0000;
        rom[9][1258] = 16'h0000;
        rom[9][1259] = 16'h0000;
        rom[9][1260] = 16'h0000;
        rom[9][1261] = 16'h0000;
        rom[9][1262] = 16'h0000;
        rom[9][1263] = 16'h0000;
        rom[9][1264] = 16'h0000;
        rom[9][1265] = 16'h0000;
        rom[9][1266] = 16'h0000;
        rom[9][1267] = 16'h0000;
        rom[9][1268] = 16'h0000;
        rom[9][1269] = 16'h0000;
        rom[9][1270] = 16'h0000;
        rom[9][1271] = 16'h0000;
        rom[9][1272] = 16'h0000;
        rom[9][1273] = 16'h0000;
    end

    always @(*) begin
        data_out = rom[addr][index];
    end
endmodule
