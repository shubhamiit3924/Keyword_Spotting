// Q8.8 Fixed-Point ROM: rom_layer2_weights
module rom_layer2_weights (
    input [7:0] addr,
    input [6:0] index,
    output reg signed [15:0] data_out
);

    reg signed [15:0] rom [0:255][0:127];

    initial begin
        rom[0][0] = 16'hFFD9;
        rom[0][1] = 16'h0011;
        rom[0][2] = 16'h0004;
        rom[0][3] = 16'h001B;
        rom[0][4] = 16'h001D;
        rom[0][5] = 16'h0029;
        rom[0][6] = 16'hFFCF;
        rom[0][7] = 16'h0002;
        rom[0][8] = 16'h0011;
        rom[0][9] = 16'h0013;
        rom[0][10] = 16'h001E;
        rom[0][11] = 16'h0017;
        rom[0][12] = 16'hFFE1;
        rom[0][13] = 16'hFFFE;
        rom[0][14] = 16'hFFEC;
        rom[0][15] = 16'h000A;
        rom[0][16] = 16'hFFC8;
        rom[0][17] = 16'hFFF8;
        rom[0][18] = 16'h0011;
        rom[0][19] = 16'h000D;
        rom[0][20] = 16'hFFED;
        rom[0][21] = 16'h0000;
        rom[0][22] = 16'hFFF6;
        rom[0][23] = 16'hFFF9;
        rom[0][24] = 16'h0015;
        rom[0][25] = 16'hFFD1;
        rom[0][26] = 16'h0007;
        rom[0][27] = 16'h0017;
        rom[0][28] = 16'h000F;
        rom[0][29] = 16'hFFFF;
        rom[0][30] = 16'hFFF7;
        rom[0][31] = 16'hFFEE;
        rom[0][32] = 16'hFFFF;
        rom[0][33] = 16'h0017;
        rom[0][34] = 16'hFFE8;
        rom[0][35] = 16'hFFE5;
        rom[0][36] = 16'hFFE6;
        rom[0][37] = 16'h0019;
        rom[0][38] = 16'h0005;
        rom[0][39] = 16'hFFEB;
        rom[0][40] = 16'hFFF8;
        rom[0][41] = 16'h001A;
        rom[0][42] = 16'hFFE2;
        rom[0][43] = 16'hFFFF;
        rom[0][44] = 16'hFFC6;
        rom[0][45] = 16'h001B;
        rom[0][46] = 16'hFFDB;
        rom[0][47] = 16'hFFFE;
        rom[0][48] = 16'h0013;
        rom[0][49] = 16'hFFBF;
        rom[0][50] = 16'hFFFE;
        rom[0][51] = 16'hFFC1;
        rom[0][52] = 16'hFFDF;
        rom[0][53] = 16'hFFEF;
        rom[0][54] = 16'hFFD1;
        rom[0][55] = 16'hFFD7;
        rom[0][56] = 16'h0008;
        rom[0][57] = 16'hFFB2;
        rom[0][58] = 16'hFFD8;
        rom[0][59] = 16'h000D;
        rom[0][60] = 16'h0006;
        rom[0][61] = 16'h001F;
        rom[0][62] = 16'hFFBD;
        rom[0][63] = 16'hFFEA;
        rom[0][64] = 16'hFFFC;
        rom[0][65] = 16'hFFDA;
        rom[0][66] = 16'h0026;
        rom[0][67] = 16'hFFF4;
        rom[0][68] = 16'hFFC9;
        rom[0][69] = 16'h0004;
        rom[0][70] = 16'h0021;
        rom[0][71] = 16'hFFDD;
        rom[0][72] = 16'hFFF9;
        rom[0][73] = 16'h001E;
        rom[0][74] = 16'hFFDC;
        rom[0][75] = 16'h0008;
        rom[0][76] = 16'h0007;
        rom[0][77] = 16'hFFF2;
        rom[0][78] = 16'hFFEF;
        rom[0][79] = 16'hFFB0;
        rom[0][80] = 16'h001B;
        rom[0][81] = 16'hFFCD;
        rom[0][82] = 16'hFFF6;
        rom[0][83] = 16'hFFE0;
        rom[0][84] = 16'hFFD2;
        rom[0][85] = 16'h000E;
        rom[0][86] = 16'h001F;
        rom[0][87] = 16'hFFD5;
        rom[0][88] = 16'hFFE5;
        rom[0][89] = 16'hFFC8;
        rom[0][90] = 16'hFFF7;
        rom[0][91] = 16'hFFC9;
        rom[0][92] = 16'h0006;
        rom[0][93] = 16'hFFF9;
        rom[0][94] = 16'hFFF4;
        rom[0][95] = 16'hFFD9;
        rom[0][96] = 16'hFFEC;
        rom[0][97] = 16'hFFA8;
        rom[0][98] = 16'hFFF6;
        rom[0][99] = 16'hFFC8;
        rom[0][100] = 16'h0013;
        rom[0][101] = 16'hFFEA;
        rom[0][102] = 16'hFFE6;
        rom[0][103] = 16'hFFD9;
        rom[0][104] = 16'hFFD4;
        rom[0][105] = 16'h001B;
        rom[0][106] = 16'h0021;
        rom[0][107] = 16'h001F;
        rom[0][108] = 16'hFFC8;
        rom[0][109] = 16'hFFF9;
        rom[0][110] = 16'h0032;
        rom[0][111] = 16'h0036;
        rom[0][112] = 16'hFFA5;
        rom[0][113] = 16'hFFC9;
        rom[0][114] = 16'h001D;
        rom[0][115] = 16'hFFC5;
        rom[0][116] = 16'h0008;
        rom[0][117] = 16'hFFF8;
        rom[0][118] = 16'hFFFE;
        rom[0][119] = 16'h001B;
        rom[0][120] = 16'hFFFC;
        rom[0][121] = 16'h0020;
        rom[0][122] = 16'hFFED;
        rom[0][123] = 16'h0006;
        rom[0][124] = 16'h0000;
        rom[0][125] = 16'hFFED;
        rom[0][126] = 16'h0017;
        rom[0][127] = 16'hFFFA;
        rom[1][0] = 16'hFFE6;
        rom[1][1] = 16'h0015;
        rom[1][2] = 16'hFFFB;
        rom[1][3] = 16'hFFC8;
        rom[1][4] = 16'h0014;
        rom[1][5] = 16'h0001;
        rom[1][6] = 16'h001E;
        rom[1][7] = 16'hFFEF;
        rom[1][8] = 16'hFFD2;
        rom[1][9] = 16'hFFC1;
        rom[1][10] = 16'hFFC2;
        rom[1][11] = 16'hFFCF;
        rom[1][12] = 16'h000A;
        rom[1][13] = 16'h0009;
        rom[1][14] = 16'hFFE7;
        rom[1][15] = 16'hFFF9;
        rom[1][16] = 16'h0016;
        rom[1][17] = 16'hFFFF;
        rom[1][18] = 16'hFFAF;
        rom[1][19] = 16'hFFBF;
        rom[1][20] = 16'hFFA6;
        rom[1][21] = 16'h0018;
        rom[1][22] = 16'hFFE8;
        rom[1][23] = 16'hFFEF;
        rom[1][24] = 16'hFFF9;
        rom[1][25] = 16'hFFE9;
        rom[1][26] = 16'h0011;
        rom[1][27] = 16'hFFF4;
        rom[1][28] = 16'hFFFA;
        rom[1][29] = 16'hFFEB;
        rom[1][30] = 16'h001A;
        rom[1][31] = 16'hFFEB;
        rom[1][32] = 16'hFFF5;
        rom[1][33] = 16'hFFBD;
        rom[1][34] = 16'hFFFD;
        rom[1][35] = 16'h000C;
        rom[1][36] = 16'h0006;
        rom[1][37] = 16'hFFD7;
        rom[1][38] = 16'hFFE5;
        rom[1][39] = 16'h001A;
        rom[1][40] = 16'hFFD9;
        rom[1][41] = 16'hFFFD;
        rom[1][42] = 16'hFFF1;
        rom[1][43] = 16'h001E;
        rom[1][44] = 16'hFFF3;
        rom[1][45] = 16'hFFF8;
        rom[1][46] = 16'hFFFE;
        rom[1][47] = 16'hFFFE;
        rom[1][48] = 16'h0022;
        rom[1][49] = 16'h0002;
        rom[1][50] = 16'hFFFB;
        rom[1][51] = 16'h001A;
        rom[1][52] = 16'hFFE2;
        rom[1][53] = 16'hFFF6;
        rom[1][54] = 16'h0023;
        rom[1][55] = 16'h0001;
        rom[1][56] = 16'h002A;
        rom[1][57] = 16'h0013;
        rom[1][58] = 16'hFFEE;
        rom[1][59] = 16'hFFC0;
        rom[1][60] = 16'h0038;
        rom[1][61] = 16'hFFE1;
        rom[1][62] = 16'h0002;
        rom[1][63] = 16'h001F;
        rom[1][64] = 16'hFFDC;
        rom[1][65] = 16'hFFDF;
        rom[1][66] = 16'h0004;
        rom[1][67] = 16'h0007;
        rom[1][68] = 16'h0000;
        rom[1][69] = 16'h000B;
        rom[1][70] = 16'h000F;
        rom[1][71] = 16'hFFE6;
        rom[1][72] = 16'h0018;
        rom[1][73] = 16'h0015;
        rom[1][74] = 16'h0002;
        rom[1][75] = 16'hFFC8;
        rom[1][76] = 16'hFFEE;
        rom[1][77] = 16'h000C;
        rom[1][78] = 16'hFFFC;
        rom[1][79] = 16'hFFF7;
        rom[1][80] = 16'h000A;
        rom[1][81] = 16'h0010;
        rom[1][82] = 16'hFFFD;
        rom[1][83] = 16'hFFED;
        rom[1][84] = 16'h0005;
        rom[1][85] = 16'h000A;
        rom[1][86] = 16'hFFDA;
        rom[1][87] = 16'hFFC4;
        rom[1][88] = 16'hFFDE;
        rom[1][89] = 16'h0014;
        rom[1][90] = 16'hFFE2;
        rom[1][91] = 16'hFFA7;
        rom[1][92] = 16'hFFD0;
        rom[1][93] = 16'hFFF5;
        rom[1][94] = 16'hFFE1;
        rom[1][95] = 16'hFFD5;
        rom[1][96] = 16'h001E;
        rom[1][97] = 16'h0015;
        rom[1][98] = 16'h0004;
        rom[1][99] = 16'hFFEF;
        rom[1][100] = 16'hFFDC;
        rom[1][101] = 16'hFFDB;
        rom[1][102] = 16'h0002;
        rom[1][103] = 16'h0027;
        rom[1][104] = 16'hFFFD;
        rom[1][105] = 16'h001A;
        rom[1][106] = 16'h000A;
        rom[1][107] = 16'hFFEC;
        rom[1][108] = 16'hFFE8;
        rom[1][109] = 16'hFFE5;
        rom[1][110] = 16'h0006;
        rom[1][111] = 16'hFFEC;
        rom[1][112] = 16'hFFE3;
        rom[1][113] = 16'h0020;
        rom[1][114] = 16'h000C;
        rom[1][115] = 16'h000A;
        rom[1][116] = 16'hFFD2;
        rom[1][117] = 16'hFFE2;
        rom[1][118] = 16'h0026;
        rom[1][119] = 16'hFFFD;
        rom[1][120] = 16'h0007;
        rom[1][121] = 16'hFFEF;
        rom[1][122] = 16'hFFDF;
        rom[1][123] = 16'hFFF9;
        rom[1][124] = 16'hFFF8;
        rom[1][125] = 16'h0011;
        rom[1][126] = 16'hFFD2;
        rom[1][127] = 16'hFFE1;
        rom[2][0] = 16'h0011;
        rom[2][1] = 16'h0000;
        rom[2][2] = 16'h0012;
        rom[2][3] = 16'hFFFC;
        rom[2][4] = 16'hFFFE;
        rom[2][5] = 16'h000F;
        rom[2][6] = 16'hFFBF;
        rom[2][7] = 16'h0007;
        rom[2][8] = 16'h0002;
        rom[2][9] = 16'hFFE8;
        rom[2][10] = 16'h000B;
        rom[2][11] = 16'h002E;
        rom[2][12] = 16'hFFE3;
        rom[2][13] = 16'hFFEC;
        rom[2][14] = 16'hFFD3;
        rom[2][15] = 16'hFFFF;
        rom[2][16] = 16'hFFBA;
        rom[2][17] = 16'h0005;
        rom[2][18] = 16'h0046;
        rom[2][19] = 16'h0012;
        rom[2][20] = 16'h0046;
        rom[2][21] = 16'hFFF8;
        rom[2][22] = 16'hFFF9;
        rom[2][23] = 16'h0039;
        rom[2][24] = 16'hFFF9;
        rom[2][25] = 16'hFFDC;
        rom[2][26] = 16'h002F;
        rom[2][27] = 16'hFFFB;
        rom[2][28] = 16'hFFE5;
        rom[2][29] = 16'hFFC1;
        rom[2][30] = 16'hFFFC;
        rom[2][31] = 16'hFFE9;
        rom[2][32] = 16'h002C;
        rom[2][33] = 16'h0011;
        rom[2][34] = 16'hFFFE;
        rom[2][35] = 16'hFFE5;
        rom[2][36] = 16'hFFFA;
        rom[2][37] = 16'hFFF7;
        rom[2][38] = 16'h0010;
        rom[2][39] = 16'hFFB4;
        rom[2][40] = 16'hFFE1;
        rom[2][41] = 16'hFFF8;
        rom[2][42] = 16'hFFD4;
        rom[2][43] = 16'h0013;
        rom[2][44] = 16'hFFE1;
        rom[2][45] = 16'h001F;
        rom[2][46] = 16'h001B;
        rom[2][47] = 16'hFFE1;
        rom[2][48] = 16'hFFFD;
        rom[2][49] = 16'hFFF9;
        rom[2][50] = 16'h000D;
        rom[2][51] = 16'hFFF7;
        rom[2][52] = 16'h0010;
        rom[2][53] = 16'h0029;
        rom[2][54] = 16'h0027;
        rom[2][55] = 16'hFFF4;
        rom[2][56] = 16'hFFEE;
        rom[2][57] = 16'h0019;
        rom[2][58] = 16'h0011;
        rom[2][59] = 16'h0020;
        rom[2][60] = 16'hFFC6;
        rom[2][61] = 16'hFFC1;
        rom[2][62] = 16'h000D;
        rom[2][63] = 16'hFFE1;
        rom[2][64] = 16'hFFE7;
        rom[2][65] = 16'hFFFE;
        rom[2][66] = 16'h0014;
        rom[2][67] = 16'h0009;
        rom[2][68] = 16'hFFCB;
        rom[2][69] = 16'hFFDD;
        rom[2][70] = 16'h0006;
        rom[2][71] = 16'hFFFB;
        rom[2][72] = 16'h0009;
        rom[2][73] = 16'h001A;
        rom[2][74] = 16'hFFB2;
        rom[2][75] = 16'hFFF6;
        rom[2][76] = 16'hFFF6;
        rom[2][77] = 16'hFFF2;
        rom[2][78] = 16'h0016;
        rom[2][79] = 16'hFFFE;
        rom[2][80] = 16'hFFED;
        rom[2][81] = 16'h0021;
        rom[2][82] = 16'h0011;
        rom[2][83] = 16'hFFE0;
        rom[2][84] = 16'hFFF1;
        rom[2][85] = 16'h0017;
        rom[2][86] = 16'hFFFC;
        rom[2][87] = 16'h000D;
        rom[2][88] = 16'hFFFD;
        rom[2][89] = 16'h0032;
        rom[2][90] = 16'h002C;
        rom[2][91] = 16'hFFFE;
        rom[2][92] = 16'h0008;
        rom[2][93] = 16'hFFF9;
        rom[2][94] = 16'hFFF3;
        rom[2][95] = 16'h001D;
        rom[2][96] = 16'h001C;
        rom[2][97] = 16'h0002;
        rom[2][98] = 16'hFFB5;
        rom[2][99] = 16'hFFFE;
        rom[2][100] = 16'hFFC7;
        rom[2][101] = 16'h0002;
        rom[2][102] = 16'hFFF2;
        rom[2][103] = 16'h0000;
        rom[2][104] = 16'h001E;
        rom[2][105] = 16'h0018;
        rom[2][106] = 16'hFFEA;
        rom[2][107] = 16'hFFFE;
        rom[2][108] = 16'h0011;
        rom[2][109] = 16'hFFEE;
        rom[2][110] = 16'h0018;
        rom[2][111] = 16'hFFFF;
        rom[2][112] = 16'hFFEE;
        rom[2][113] = 16'hFFBD;
        rom[2][114] = 16'hFFCB;
        rom[2][115] = 16'hFFEE;
        rom[2][116] = 16'h001E;
        rom[2][117] = 16'hFFDF;
        rom[2][118] = 16'h001A;
        rom[2][119] = 16'h0006;
        rom[2][120] = 16'h0005;
        rom[2][121] = 16'hFFFA;
        rom[2][122] = 16'h0033;
        rom[2][123] = 16'h002A;
        rom[2][124] = 16'h0019;
        rom[2][125] = 16'h0017;
        rom[2][126] = 16'h0029;
        rom[2][127] = 16'h0001;
        rom[3][0] = 16'hFFEB;
        rom[3][1] = 16'hFFEC;
        rom[3][2] = 16'hFFF4;
        rom[3][3] = 16'hFFC9;
        rom[3][4] = 16'hFFBA;
        rom[3][5] = 16'hFFF2;
        rom[3][6] = 16'h001A;
        rom[3][7] = 16'h001B;
        rom[3][8] = 16'hFFED;
        rom[3][9] = 16'hFFDD;
        rom[3][10] = 16'hFFBA;
        rom[3][11] = 16'h000E;
        rom[3][12] = 16'h001B;
        rom[3][13] = 16'hFFF8;
        rom[3][14] = 16'hFFE5;
        rom[3][15] = 16'h000C;
        rom[3][16] = 16'h000D;
        rom[3][17] = 16'hFFF5;
        rom[3][18] = 16'hFFFC;
        rom[3][19] = 16'hFFEF;
        rom[3][20] = 16'hFFD4;
        rom[3][21] = 16'h0020;
        rom[3][22] = 16'h0010;
        rom[3][23] = 16'hFFFD;
        rom[3][24] = 16'h0008;
        rom[3][25] = 16'h000A;
        rom[3][26] = 16'hFFF0;
        rom[3][27] = 16'hFFF5;
        rom[3][28] = 16'h0016;
        rom[3][29] = 16'h0034;
        rom[3][30] = 16'h001D;
        rom[3][31] = 16'h000C;
        rom[3][32] = 16'hFFE5;
        rom[3][33] = 16'h001A;
        rom[3][34] = 16'h0007;
        rom[3][35] = 16'h001B;
        rom[3][36] = 16'h0017;
        rom[3][37] = 16'hFFE5;
        rom[3][38] = 16'hFFF1;
        rom[3][39] = 16'h001F;
        rom[3][40] = 16'h001B;
        rom[3][41] = 16'hFFE2;
        rom[3][42] = 16'h0004;
        rom[3][43] = 16'hFFBE;
        rom[3][44] = 16'h0005;
        rom[3][45] = 16'h0008;
        rom[3][46] = 16'hFFF4;
        rom[3][47] = 16'h0008;
        rom[3][48] = 16'h000F;
        rom[3][49] = 16'h0005;
        rom[3][50] = 16'h0003;
        rom[3][51] = 16'hFFE4;
        rom[3][52] = 16'h0016;
        rom[3][53] = 16'h001C;
        rom[3][54] = 16'h0011;
        rom[3][55] = 16'h0016;
        rom[3][56] = 16'hFFDC;
        rom[3][57] = 16'hFFBE;
        rom[3][58] = 16'h000B;
        rom[3][59] = 16'hFFE1;
        rom[3][60] = 16'hFFFE;
        rom[3][61] = 16'h001A;
        rom[3][62] = 16'h0027;
        rom[3][63] = 16'h0014;
        rom[3][64] = 16'hFFC8;
        rom[3][65] = 16'h001A;
        rom[3][66] = 16'hFFF0;
        rom[3][67] = 16'hFFE1;
        rom[3][68] = 16'h001C;
        rom[3][69] = 16'hFFF2;
        rom[3][70] = 16'h000F;
        rom[3][71] = 16'hFFF4;
        rom[3][72] = 16'h000E;
        rom[3][73] = 16'hFFF3;
        rom[3][74] = 16'h0018;
        rom[3][75] = 16'h000C;
        rom[3][76] = 16'hFFF5;
        rom[3][77] = 16'hFFE7;
        rom[3][78] = 16'hFFE5;
        rom[3][79] = 16'hFFED;
        rom[3][80] = 16'h0009;
        rom[3][81] = 16'h001E;
        rom[3][82] = 16'hFFCB;
        rom[3][83] = 16'h0007;
        rom[3][84] = 16'hFFF4;
        rom[3][85] = 16'hFFBA;
        rom[3][86] = 16'hFFC7;
        rom[3][87] = 16'hFFC1;
        rom[3][88] = 16'hFFDF;
        rom[3][89] = 16'h0007;
        rom[3][90] = 16'hFFB9;
        rom[3][91] = 16'h0000;
        rom[3][92] = 16'h0015;
        rom[3][93] = 16'h0026;
        rom[3][94] = 16'h000E;
        rom[3][95] = 16'hFFBD;
        rom[3][96] = 16'hFFF5;
        rom[3][97] = 16'h0003;
        rom[3][98] = 16'h0000;
        rom[3][99] = 16'h000E;
        rom[3][100] = 16'hFFFA;
        rom[3][101] = 16'hFFDC;
        rom[3][102] = 16'h0009;
        rom[3][103] = 16'hFFB0;
        rom[3][104] = 16'hFFC6;
        rom[3][105] = 16'hFFC6;
        rom[3][106] = 16'hFFF1;
        rom[3][107] = 16'h0002;
        rom[3][108] = 16'hFFFF;
        rom[3][109] = 16'h000A;
        rom[3][110] = 16'hFFE9;
        rom[3][111] = 16'h000F;
        rom[3][112] = 16'hFFE2;
        rom[3][113] = 16'hFFE1;
        rom[3][114] = 16'hFFFE;
        rom[3][115] = 16'hFFFB;
        rom[3][116] = 16'hFFFD;
        rom[3][117] = 16'hFFC3;
        rom[3][118] = 16'hFFDE;
        rom[3][119] = 16'h0038;
        rom[3][120] = 16'h000B;
        rom[3][121] = 16'hFFCB;
        rom[3][122] = 16'h0010;
        rom[3][123] = 16'h0002;
        rom[3][124] = 16'hFFF7;
        rom[3][125] = 16'hFFDA;
        rom[3][126] = 16'hFFEF;
        rom[3][127] = 16'hFFFE;
        rom[4][0] = 16'hFFC6;
        rom[4][1] = 16'h0018;
        rom[4][2] = 16'h001A;
        rom[4][3] = 16'hFFF4;
        rom[4][4] = 16'h0017;
        rom[4][5] = 16'h0034;
        rom[4][6] = 16'hFFF2;
        rom[4][7] = 16'h0011;
        rom[4][8] = 16'hFFEB;
        rom[4][9] = 16'h0013;
        rom[4][10] = 16'hFFE5;
        rom[4][11] = 16'hFFED;
        rom[4][12] = 16'hFFF9;
        rom[4][13] = 16'h0001;
        rom[4][14] = 16'h000B;
        rom[4][15] = 16'h001F;
        rom[4][16] = 16'hFFE0;
        rom[4][17] = 16'h000A;
        rom[4][18] = 16'hFFF9;
        rom[4][19] = 16'h0001;
        rom[4][20] = 16'hFFEF;
        rom[4][21] = 16'h0015;
        rom[4][22] = 16'h0011;
        rom[4][23] = 16'hFFF4;
        rom[4][24] = 16'h0015;
        rom[4][25] = 16'h0016;
        rom[4][26] = 16'hFFFA;
        rom[4][27] = 16'hFFFB;
        rom[4][28] = 16'hFFD6;
        rom[4][29] = 16'h000C;
        rom[4][30] = 16'h0024;
        rom[4][31] = 16'hFFC2;
        rom[4][32] = 16'h0015;
        rom[4][33] = 16'h0002;
        rom[4][34] = 16'hFFEA;
        rom[4][35] = 16'hFFD2;
        rom[4][36] = 16'h0010;
        rom[4][37] = 16'hFFFB;
        rom[4][38] = 16'h0025;
        rom[4][39] = 16'hFFE1;
        rom[4][40] = 16'hFFB0;
        rom[4][41] = 16'hFFF4;
        rom[4][42] = 16'h0004;
        rom[4][43] = 16'hFFDC;
        rom[4][44] = 16'hFFDE;
        rom[4][45] = 16'hFFD1;
        rom[4][46] = 16'h0007;
        rom[4][47] = 16'h0002;
        rom[4][48] = 16'hFFEF;
        rom[4][49] = 16'h001F;
        rom[4][50] = 16'h001D;
        rom[4][51] = 16'hFFE4;
        rom[4][52] = 16'hFFDE;
        rom[4][53] = 16'hFFD9;
        rom[4][54] = 16'hFFD7;
        rom[4][55] = 16'hFFE1;
        rom[4][56] = 16'h0021;
        rom[4][57] = 16'hFFD3;
        rom[4][58] = 16'hFFF8;
        rom[4][59] = 16'hFFD0;
        rom[4][60] = 16'h0024;
        rom[4][61] = 16'h001B;
        rom[4][62] = 16'h0000;
        rom[4][63] = 16'h000F;
        rom[4][64] = 16'h0013;
        rom[4][65] = 16'hFFE4;
        rom[4][66] = 16'h0016;
        rom[4][67] = 16'h0027;
        rom[4][68] = 16'hFFDF;
        rom[4][69] = 16'h0008;
        rom[4][70] = 16'h001C;
        rom[4][71] = 16'hFFDD;
        rom[4][72] = 16'hFFD2;
        rom[4][73] = 16'h0011;
        rom[4][74] = 16'hFFDC;
        rom[4][75] = 16'h001F;
        rom[4][76] = 16'h001B;
        rom[4][77] = 16'hFFFF;
        rom[4][78] = 16'h0010;
        rom[4][79] = 16'hFFF4;
        rom[4][80] = 16'h0000;
        rom[4][81] = 16'hFFD5;
        rom[4][82] = 16'h000D;
        rom[4][83] = 16'hFFFE;
        rom[4][84] = 16'h0008;
        rom[4][85] = 16'h0019;
        rom[4][86] = 16'hFFCB;
        rom[4][87] = 16'h000E;
        rom[4][88] = 16'hFFE7;
        rom[4][89] = 16'hFFF5;
        rom[4][90] = 16'h000C;
        rom[4][91] = 16'hFFCD;
        rom[4][92] = 16'h0004;
        rom[4][93] = 16'hFFAB;
        rom[4][94] = 16'hFFAD;
        rom[4][95] = 16'hFFCA;
        rom[4][96] = 16'hFFF9;
        rom[4][97] = 16'hFFD9;
        rom[4][98] = 16'hFFDC;
        rom[4][99] = 16'hFFF6;
        rom[4][100] = 16'hFFDC;
        rom[4][101] = 16'hFFE5;
        rom[4][102] = 16'hFFE6;
        rom[4][103] = 16'hFFE3;
        rom[4][104] = 16'hFFE1;
        rom[4][105] = 16'hFFC2;
        rom[4][106] = 16'h0028;
        rom[4][107] = 16'hFFDF;
        rom[4][108] = 16'hFFEA;
        rom[4][109] = 16'hFFEF;
        rom[4][110] = 16'h001A;
        rom[4][111] = 16'hFFEA;
        rom[4][112] = 16'hFFFB;
        rom[4][113] = 16'hFFF6;
        rom[4][114] = 16'hFFDC;
        rom[4][115] = 16'hFFAF;
        rom[4][116] = 16'h0004;
        rom[4][117] = 16'h0033;
        rom[4][118] = 16'h002D;
        rom[4][119] = 16'h000F;
        rom[4][120] = 16'h0001;
        rom[4][121] = 16'hFFF2;
        rom[4][122] = 16'hFFE7;
        rom[4][123] = 16'hFFFC;
        rom[4][124] = 16'hFFEE;
        rom[4][125] = 16'hFFF4;
        rom[4][126] = 16'hFFB3;
        rom[4][127] = 16'hFFF6;
        rom[5][0] = 16'h0008;
        rom[5][1] = 16'h0003;
        rom[5][2] = 16'hFFD2;
        rom[5][3] = 16'hFFF9;
        rom[5][4] = 16'hFFDD;
        rom[5][5] = 16'hFFFE;
        rom[5][6] = 16'hFFDA;
        rom[5][7] = 16'h0002;
        rom[5][8] = 16'hFFBC;
        rom[5][9] = 16'h000F;
        rom[5][10] = 16'h000E;
        rom[5][11] = 16'h0001;
        rom[5][12] = 16'h0011;
        rom[5][13] = 16'h0008;
        rom[5][14] = 16'hFFBE;
        rom[5][15] = 16'hFFF4;
        rom[5][16] = 16'hFFDC;
        rom[5][17] = 16'hFFFC;
        rom[5][18] = 16'hFFEE;
        rom[5][19] = 16'hFFE4;
        rom[5][20] = 16'h0028;
        rom[5][21] = 16'hFFED;
        rom[5][22] = 16'hFFEF;
        rom[5][23] = 16'h000A;
        rom[5][24] = 16'hFFFF;
        rom[5][25] = 16'hFFE5;
        rom[5][26] = 16'h000E;
        rom[5][27] = 16'hFFFB;
        rom[5][28] = 16'h0025;
        rom[5][29] = 16'h0003;
        rom[5][30] = 16'hFFFE;
        rom[5][31] = 16'hFFD4;
        rom[5][32] = 16'hFFFE;
        rom[5][33] = 16'h0015;
        rom[5][34] = 16'hFFE5;
        rom[5][35] = 16'hFFE1;
        rom[5][36] = 16'h0009;
        rom[5][37] = 16'hFFF4;
        rom[5][38] = 16'h001E;
        rom[5][39] = 16'hFFDC;
        rom[5][40] = 16'hFFF8;
        rom[5][41] = 16'h000A;
        rom[5][42] = 16'h002C;
        rom[5][43] = 16'h0020;
        rom[5][44] = 16'hFFF4;
        rom[5][45] = 16'hFFDA;
        rom[5][46] = 16'h000F;
        rom[5][47] = 16'hFFDC;
        rom[5][48] = 16'h0008;
        rom[5][49] = 16'h0021;
        rom[5][50] = 16'hFFEC;
        rom[5][51] = 16'h0006;
        rom[5][52] = 16'hFFE5;
        rom[5][53] = 16'hFFFD;
        rom[5][54] = 16'hFFC2;
        rom[5][55] = 16'h0006;
        rom[5][56] = 16'h0007;
        rom[5][57] = 16'h0009;
        rom[5][58] = 16'hFFF7;
        rom[5][59] = 16'h0024;
        rom[5][60] = 16'hFFE1;
        rom[5][61] = 16'h005A;
        rom[5][62] = 16'hFFD4;
        rom[5][63] = 16'h000F;
        rom[5][64] = 16'h0021;
        rom[5][65] = 16'hFFC4;
        rom[5][66] = 16'hFFFF;
        rom[5][67] = 16'h0032;
        rom[5][68] = 16'hFFEE;
        rom[5][69] = 16'h0010;
        rom[5][70] = 16'hFFFE;
        rom[5][71] = 16'hFFD0;
        rom[5][72] = 16'hFFFC;
        rom[5][73] = 16'h0004;
        rom[5][74] = 16'hFFC3;
        rom[5][75] = 16'hFFFE;
        rom[5][76] = 16'h0018;
        rom[5][77] = 16'h0003;
        rom[5][78] = 16'hFFFF;
        rom[5][79] = 16'h001B;
        rom[5][80] = 16'h000C;
        rom[5][81] = 16'hFFF4;
        rom[5][82] = 16'h002E;
        rom[5][83] = 16'hFFEE;
        rom[5][84] = 16'h001E;
        rom[5][85] = 16'h0018;
        rom[5][86] = 16'hFFF9;
        rom[5][87] = 16'h0002;
        rom[5][88] = 16'hFFCB;
        rom[5][89] = 16'hFFC6;
        rom[5][90] = 16'h0011;
        rom[5][91] = 16'hFFEF;
        rom[5][92] = 16'hFFE5;
        rom[5][93] = 16'hFFE6;
        rom[5][94] = 16'h0026;
        rom[5][95] = 16'hFFE5;
        rom[5][96] = 16'hFFE9;
        rom[5][97] = 16'h001C;
        rom[5][98] = 16'hFFF4;
        rom[5][99] = 16'h0028;
        rom[5][100] = 16'hFFFC;
        rom[5][101] = 16'hFFF4;
        rom[5][102] = 16'hFFF3;
        rom[5][103] = 16'h0010;
        rom[5][104] = 16'h0006;
        rom[5][105] = 16'hFFDC;
        rom[5][106] = 16'hFFED;
        rom[5][107] = 16'h0006;
        rom[5][108] = 16'h0000;
        rom[5][109] = 16'hFFF0;
        rom[5][110] = 16'h001E;
        rom[5][111] = 16'h0020;
        rom[5][112] = 16'h0019;
        rom[5][113] = 16'hFFD2;
        rom[5][114] = 16'h000C;
        rom[5][115] = 16'hFFFE;
        rom[5][116] = 16'hFFFA;
        rom[5][117] = 16'hFFF1;
        rom[5][118] = 16'hFFF0;
        rom[5][119] = 16'h0024;
        rom[5][120] = 16'h0003;
        rom[5][121] = 16'h0017;
        rom[5][122] = 16'h0007;
        rom[5][123] = 16'hFFE6;
        rom[5][124] = 16'hFFC7;
        rom[5][125] = 16'hFFF5;
        rom[5][126] = 16'hFFD9;
        rom[5][127] = 16'h0005;
        rom[6][0] = 16'hFFFD;
        rom[6][1] = 16'h0025;
        rom[6][2] = 16'h001B;
        rom[6][3] = 16'hFFD2;
        rom[6][4] = 16'h0019;
        rom[6][5] = 16'h0009;
        rom[6][6] = 16'h0021;
        rom[6][7] = 16'h0005;
        rom[6][8] = 16'h0007;
        rom[6][9] = 16'hFFFD;
        rom[6][10] = 16'hFFD2;
        rom[6][11] = 16'hFFE6;
        rom[6][12] = 16'hFFCD;
        rom[6][13] = 16'h0011;
        rom[6][14] = 16'hFFEE;
        rom[6][15] = 16'hFFDB;
        rom[6][16] = 16'h002C;
        rom[6][17] = 16'hFFC6;
        rom[6][18] = 16'h0024;
        rom[6][19] = 16'hFFFE;
        rom[6][20] = 16'hFFED;
        rom[6][21] = 16'h0014;
        rom[6][22] = 16'h0016;
        rom[6][23] = 16'h0003;
        rom[6][24] = 16'hFFB6;
        rom[6][25] = 16'h002C;
        rom[6][26] = 16'hFFF6;
        rom[6][27] = 16'hFFEF;
        rom[6][28] = 16'hFFDB;
        rom[6][29] = 16'h0006;
        rom[6][30] = 16'h0029;
        rom[6][31] = 16'hFFCF;
        rom[6][32] = 16'h0019;
        rom[6][33] = 16'hFFCD;
        rom[6][34] = 16'h0013;
        rom[6][35] = 16'hFFD7;
        rom[6][36] = 16'h0026;
        rom[6][37] = 16'hFFC7;
        rom[6][38] = 16'hFFC2;
        rom[6][39] = 16'h000C;
        rom[6][40] = 16'h0021;
        rom[6][41] = 16'h002F;
        rom[6][42] = 16'hFFEA;
        rom[6][43] = 16'h0007;
        rom[6][44] = 16'h001D;
        rom[6][45] = 16'hFFC4;
        rom[6][46] = 16'h001E;
        rom[6][47] = 16'h000B;
        rom[6][48] = 16'h0003;
        rom[6][49] = 16'hFFF8;
        rom[6][50] = 16'hFFFA;
        rom[6][51] = 16'hFFF3;
        rom[6][52] = 16'hFFFC;
        rom[6][53] = 16'hFFF9;
        rom[6][54] = 16'h0012;
        rom[6][55] = 16'h0009;
        rom[6][56] = 16'hFFE3;
        rom[6][57] = 16'h0019;
        rom[6][58] = 16'hFFDC;
        rom[6][59] = 16'hFFCA;
        rom[6][60] = 16'hFFEB;
        rom[6][61] = 16'hFFD7;
        rom[6][62] = 16'h000E;
        rom[6][63] = 16'h0013;
        rom[6][64] = 16'h0026;
        rom[6][65] = 16'hFFF8;
        rom[6][66] = 16'h001A;
        rom[6][67] = 16'h000C;
        rom[6][68] = 16'hFFD7;
        rom[6][69] = 16'h0019;
        rom[6][70] = 16'hFFBA;
        rom[6][71] = 16'h001C;
        rom[6][72] = 16'hFFBA;
        rom[6][73] = 16'hFFFB;
        rom[6][74] = 16'hFFB4;
        rom[6][75] = 16'hFFCA;
        rom[6][76] = 16'hFFFC;
        rom[6][77] = 16'hFFCD;
        rom[6][78] = 16'h0002;
        rom[6][79] = 16'h0016;
        rom[6][80] = 16'hFFF8;
        rom[6][81] = 16'h000A;
        rom[6][82] = 16'h000F;
        rom[6][83] = 16'h001F;
        rom[6][84] = 16'hFFE5;
        rom[6][85] = 16'hFFD9;
        rom[6][86] = 16'hFFDE;
        rom[6][87] = 16'h0002;
        rom[6][88] = 16'h0017;
        rom[6][89] = 16'hFFCC;
        rom[6][90] = 16'h0002;
        rom[6][91] = 16'hFFFD;
        rom[6][92] = 16'hFFAC;
        rom[6][93] = 16'hFFDF;
        rom[6][94] = 16'h0038;
        rom[6][95] = 16'hFFF4;
        rom[6][96] = 16'h0005;
        rom[6][97] = 16'hFFF4;
        rom[6][98] = 16'hFFF9;
        rom[6][99] = 16'hFFED;
        rom[6][100] = 16'hFFFC;
        rom[6][101] = 16'h0011;
        rom[6][102] = 16'h0038;
        rom[6][103] = 16'h001B;
        rom[6][104] = 16'hFFEF;
        rom[6][105] = 16'h001C;
        rom[6][106] = 16'hFFF4;
        rom[6][107] = 16'hFFBD;
        rom[6][108] = 16'h0000;
        rom[6][109] = 16'hFFCB;
        rom[6][110] = 16'h0017;
        rom[6][111] = 16'hFFF7;
        rom[6][112] = 16'hFFF6;
        rom[6][113] = 16'h002B;
        rom[6][114] = 16'hFFFD;
        rom[6][115] = 16'hFFF8;
        rom[6][116] = 16'h001B;
        rom[6][117] = 16'hFFED;
        rom[6][118] = 16'hFFF1;
        rom[6][119] = 16'hFFEF;
        rom[6][120] = 16'hFFE0;
        rom[6][121] = 16'hFFC8;
        rom[6][122] = 16'hFFE1;
        rom[6][123] = 16'hFFB6;
        rom[6][124] = 16'hFFEE;
        rom[6][125] = 16'hFFDB;
        rom[6][126] = 16'hFFBA;
        rom[6][127] = 16'h0024;
        rom[7][0] = 16'h001C;
        rom[7][1] = 16'hFFD2;
        rom[7][2] = 16'h000D;
        rom[7][3] = 16'hFFD5;
        rom[7][4] = 16'hFFEA;
        rom[7][5] = 16'hFFD0;
        rom[7][6] = 16'hFFCC;
        rom[7][7] = 16'h000C;
        rom[7][8] = 16'h0029;
        rom[7][9] = 16'h0002;
        rom[7][10] = 16'hFFC7;
        rom[7][11] = 16'h0012;
        rom[7][12] = 16'hFFEA;
        rom[7][13] = 16'h0027;
        rom[7][14] = 16'hFFFF;
        rom[7][15] = 16'h0018;
        rom[7][16] = 16'hFFF0;
        rom[7][17] = 16'hFFC7;
        rom[7][18] = 16'h001F;
        rom[7][19] = 16'hFFD7;
        rom[7][20] = 16'h0012;
        rom[7][21] = 16'h0010;
        rom[7][22] = 16'hFFE6;
        rom[7][23] = 16'hFFF4;
        rom[7][24] = 16'h000E;
        rom[7][25] = 16'hFFCC;
        rom[7][26] = 16'h000F;
        rom[7][27] = 16'h0009;
        rom[7][28] = 16'hFFC6;
        rom[7][29] = 16'hFFFE;
        rom[7][30] = 16'h0030;
        rom[7][31] = 16'h0029;
        rom[7][32] = 16'hFFF9;
        rom[7][33] = 16'hFFFE;
        rom[7][34] = 16'h003D;
        rom[7][35] = 16'h0001;
        rom[7][36] = 16'h0021;
        rom[7][37] = 16'h0017;
        rom[7][38] = 16'h001F;
        rom[7][39] = 16'hFFCD;
        rom[7][40] = 16'hFFC8;
        rom[7][41] = 16'h003A;
        rom[7][42] = 16'h0019;
        rom[7][43] = 16'hFFFE;
        rom[7][44] = 16'hFFFB;
        rom[7][45] = 16'hFFE5;
        rom[7][46] = 16'h0000;
        rom[7][47] = 16'hFFC1;
        rom[7][48] = 16'hFFE1;
        rom[7][49] = 16'hFFC8;
        rom[7][50] = 16'h0001;
        rom[7][51] = 16'hFFDF;
        rom[7][52] = 16'h0006;
        rom[7][53] = 16'hFFE9;
        rom[7][54] = 16'hFFAC;
        rom[7][55] = 16'hFFC1;
        rom[7][56] = 16'h0029;
        rom[7][57] = 16'h0007;
        rom[7][58] = 16'hFFE1;
        rom[7][59] = 16'h0025;
        rom[7][60] = 16'h0009;
        rom[7][61] = 16'hFFE1;
        rom[7][62] = 16'hFFD8;
        rom[7][63] = 16'hFFCE;
        rom[7][64] = 16'h000F;
        rom[7][65] = 16'h0024;
        rom[7][66] = 16'hFFFF;
        rom[7][67] = 16'h0006;
        rom[7][68] = 16'hFFC8;
        rom[7][69] = 16'hFFC9;
        rom[7][70] = 16'h0011;
        rom[7][71] = 16'h0011;
        rom[7][72] = 16'h0024;
        rom[7][73] = 16'hFFE5;
        rom[7][74] = 16'h0028;
        rom[7][75] = 16'hFFF6;
        rom[7][76] = 16'h0026;
        rom[7][77] = 16'hFFF3;
        rom[7][78] = 16'hFFC1;
        rom[7][79] = 16'hFFFF;
        rom[7][80] = 16'hFFE8;
        rom[7][81] = 16'h0011;
        rom[7][82] = 16'hFFE1;
        rom[7][83] = 16'h0004;
        rom[7][84] = 16'h001D;
        rom[7][85] = 16'hFFD4;
        rom[7][86] = 16'h001A;
        rom[7][87] = 16'h001B;
        rom[7][88] = 16'hFFC9;
        rom[7][89] = 16'hFFB4;
        rom[7][90] = 16'hFFE2;
        rom[7][91] = 16'h001A;
        rom[7][92] = 16'hFFEF;
        rom[7][93] = 16'hFFE9;
        rom[7][94] = 16'hFFEE;
        rom[7][95] = 16'h000A;
        rom[7][96] = 16'hFFBC;
        rom[7][97] = 16'hFFE0;
        rom[7][98] = 16'hFFD0;
        rom[7][99] = 16'h001E;
        rom[7][100] = 16'hFFCF;
        rom[7][101] = 16'h0003;
        rom[7][102] = 16'h0023;
        rom[7][103] = 16'h0007;
        rom[7][104] = 16'hFFD4;
        rom[7][105] = 16'hFFE9;
        rom[7][106] = 16'h001B;
        rom[7][107] = 16'h000C;
        rom[7][108] = 16'h000B;
        rom[7][109] = 16'hFFFE;
        rom[7][110] = 16'hFFE1;
        rom[7][111] = 16'hFFED;
        rom[7][112] = 16'hFFFC;
        rom[7][113] = 16'hFFC5;
        rom[7][114] = 16'h001F;
        rom[7][115] = 16'hFFDB;
        rom[7][116] = 16'h0026;
        rom[7][117] = 16'hFFEF;
        rom[7][118] = 16'hFFD2;
        rom[7][119] = 16'hFFFB;
        rom[7][120] = 16'h0011;
        rom[7][121] = 16'hFFE9;
        rom[7][122] = 16'h0016;
        rom[7][123] = 16'h003D;
        rom[7][124] = 16'h0001;
        rom[7][125] = 16'hFFF6;
        rom[7][126] = 16'h000F;
        rom[7][127] = 16'h0000;
        rom[8][0] = 16'h000B;
        rom[8][1] = 16'h003A;
        rom[8][2] = 16'hFFE4;
        rom[8][3] = 16'hFFEF;
        rom[8][4] = 16'h002C;
        rom[8][5] = 16'hFFD2;
        rom[8][6] = 16'hFFEC;
        rom[8][7] = 16'h002F;
        rom[8][8] = 16'h000B;
        rom[8][9] = 16'h000C;
        rom[8][10] = 16'hFFEA;
        rom[8][11] = 16'hFFFB;
        rom[8][12] = 16'hFFE8;
        rom[8][13] = 16'hFFFE;
        rom[8][14] = 16'hFFCA;
        rom[8][15] = 16'h001B;
        rom[8][16] = 16'h000C;
        rom[8][17] = 16'h000B;
        rom[8][18] = 16'h000F;
        rom[8][19] = 16'h0008;
        rom[8][20] = 16'hFFE5;
        rom[8][21] = 16'hFFDA;
        rom[8][22] = 16'h0002;
        rom[8][23] = 16'h000E;
        rom[8][24] = 16'hFFF5;
        rom[8][25] = 16'hFFF1;
        rom[8][26] = 16'h0025;
        rom[8][27] = 16'hFFE7;
        rom[8][28] = 16'h0016;
        rom[8][29] = 16'h000C;
        rom[8][30] = 16'h000C;
        rom[8][31] = 16'hFFCD;
        rom[8][32] = 16'hFFC3;
        rom[8][33] = 16'hFFF9;
        rom[8][34] = 16'h0012;
        rom[8][35] = 16'hFFBC;
        rom[8][36] = 16'h0030;
        rom[8][37] = 16'h001F;
        rom[8][38] = 16'hFFF0;
        rom[8][39] = 16'hFFF3;
        rom[8][40] = 16'h0002;
        rom[8][41] = 16'hFFFC;
        rom[8][42] = 16'hFFD0;
        rom[8][43] = 16'hFFFA;
        rom[8][44] = 16'h0000;
        rom[8][45] = 16'hFFBF;
        rom[8][46] = 16'h0026;
        rom[8][47] = 16'h000C;
        rom[8][48] = 16'hFFB0;
        rom[8][49] = 16'hFFCE;
        rom[8][50] = 16'h0009;
        rom[8][51] = 16'hFFD7;
        rom[8][52] = 16'h0017;
        rom[8][53] = 16'hFFED;
        rom[8][54] = 16'hFFFB;
        rom[8][55] = 16'hFFD0;
        rom[8][56] = 16'hFFFB;
        rom[8][57] = 16'h000F;
        rom[8][58] = 16'hFFFB;
        rom[8][59] = 16'hFFEB;
        rom[8][60] = 16'h0018;
        rom[8][61] = 16'hFFDB;
        rom[8][62] = 16'hFFC4;
        rom[8][63] = 16'h0023;
        rom[8][64] = 16'hFFFA;
        rom[8][65] = 16'h0029;
        rom[8][66] = 16'hFFE6;
        rom[8][67] = 16'hFFFF;
        rom[8][68] = 16'hFFE7;
        rom[8][69] = 16'hFFDC;
        rom[8][70] = 16'hFFD9;
        rom[8][71] = 16'hFFF5;
        rom[8][72] = 16'hFFEE;
        rom[8][73] = 16'h0007;
        rom[8][74] = 16'hFFF2;
        rom[8][75] = 16'hFFFF;
        rom[8][76] = 16'hFFDF;
        rom[8][77] = 16'h0009;
        rom[8][78] = 16'hFFEB;
        rom[8][79] = 16'hFFE1;
        rom[8][80] = 16'hFFF0;
        rom[8][81] = 16'hFFDB;
        rom[8][82] = 16'hFFF4;
        rom[8][83] = 16'hFFEA;
        rom[8][84] = 16'hFFF0;
        rom[8][85] = 16'h0023;
        rom[8][86] = 16'h000D;
        rom[8][87] = 16'h0016;
        rom[8][88] = 16'hFFFE;
        rom[8][89] = 16'hFFCE;
        rom[8][90] = 16'h0010;
        rom[8][91] = 16'hFFF8;
        rom[8][92] = 16'h0003;
        rom[8][93] = 16'hFFF6;
        rom[8][94] = 16'h0035;
        rom[8][95] = 16'h0017;
        rom[8][96] = 16'hFFE2;
        rom[8][97] = 16'hFFC3;
        rom[8][98] = 16'hFFEA;
        rom[8][99] = 16'hFFED;
        rom[8][100] = 16'hFFFF;
        rom[8][101] = 16'h001F;
        rom[8][102] = 16'hFFC3;
        rom[8][103] = 16'h000C;
        rom[8][104] = 16'h0011;
        rom[8][105] = 16'h000B;
        rom[8][106] = 16'h0001;
        rom[8][107] = 16'hFFB2;
        rom[8][108] = 16'hFFAB;
        rom[8][109] = 16'hFFEC;
        rom[8][110] = 16'h0001;
        rom[8][111] = 16'hFFF8;
        rom[8][112] = 16'hFFFE;
        rom[8][113] = 16'hFFEB;
        rom[8][114] = 16'hFFE4;
        rom[8][115] = 16'h000E;
        rom[8][116] = 16'h001B;
        rom[8][117] = 16'h0019;
        rom[8][118] = 16'h0005;
        rom[8][119] = 16'hFFD4;
        rom[8][120] = 16'hFFF2;
        rom[8][121] = 16'h0019;
        rom[8][122] = 16'hFFE1;
        rom[8][123] = 16'h0012;
        rom[8][124] = 16'hFFF4;
        rom[8][125] = 16'hFFF0;
        rom[8][126] = 16'hFFD9;
        rom[8][127] = 16'h000C;
        rom[9][0] = 16'hFFEF;
        rom[9][1] = 16'h0018;
        rom[9][2] = 16'hFFEC;
        rom[9][3] = 16'hFFD6;
        rom[9][4] = 16'h0022;
        rom[9][5] = 16'hFFE4;
        rom[9][6] = 16'h0013;
        rom[9][7] = 16'h0015;
        rom[9][8] = 16'h003C;
        rom[9][9] = 16'hFFD9;
        rom[9][10] = 16'hFFD2;
        rom[9][11] = 16'h0006;
        rom[9][12] = 16'h0018;
        rom[9][13] = 16'hFFF2;
        rom[9][14] = 16'h0007;
        rom[9][15] = 16'hFFEF;
        rom[9][16] = 16'hFFFB;
        rom[9][17] = 16'h001A;
        rom[9][18] = 16'hFFD5;
        rom[9][19] = 16'h0015;
        rom[9][20] = 16'hFFF4;
        rom[9][21] = 16'hFFFD;
        rom[9][22] = 16'hFFE4;
        rom[9][23] = 16'h0026;
        rom[9][24] = 16'hFFE7;
        rom[9][25] = 16'h001D;
        rom[9][26] = 16'h000B;
        rom[9][27] = 16'hFFF9;
        rom[9][28] = 16'hFFAF;
        rom[9][29] = 16'hFFF3;
        rom[9][30] = 16'hFFEA;
        rom[9][31] = 16'hFFEB;
        rom[9][32] = 16'h0000;
        rom[9][33] = 16'hFFE9;
        rom[9][34] = 16'h000D;
        rom[9][35] = 16'hFFDA;
        rom[9][36] = 16'hFFF9;
        rom[9][37] = 16'h001E;
        rom[9][38] = 16'hFFF3;
        rom[9][39] = 16'hFFC2;
        rom[9][40] = 16'hFFEB;
        rom[9][41] = 16'h0004;
        rom[9][42] = 16'hFFDB;
        rom[9][43] = 16'h000C;
        rom[9][44] = 16'hFFD5;
        rom[9][45] = 16'hFFFC;
        rom[9][46] = 16'hFFFC;
        rom[9][47] = 16'h0006;
        rom[9][48] = 16'h0025;
        rom[9][49] = 16'h0044;
        rom[9][50] = 16'hFFF0;
        rom[9][51] = 16'hFFD0;
        rom[9][52] = 16'hFFF9;
        rom[9][53] = 16'hFFB0;
        rom[9][54] = 16'h000E;
        rom[9][55] = 16'h0014;
        rom[9][56] = 16'h0002;
        rom[9][57] = 16'hFFFC;
        rom[9][58] = 16'hFFEA;
        rom[9][59] = 16'h0044;
        rom[9][60] = 16'h0006;
        rom[9][61] = 16'hFFBB;
        rom[9][62] = 16'h0027;
        rom[9][63] = 16'h001C;
        rom[9][64] = 16'hFFF9;
        rom[9][65] = 16'h0003;
        rom[9][66] = 16'h0001;
        rom[9][67] = 16'h0004;
        rom[9][68] = 16'hFFE5;
        rom[9][69] = 16'h0007;
        rom[9][70] = 16'hFFE5;
        rom[9][71] = 16'h0009;
        rom[9][72] = 16'h002D;
        rom[9][73] = 16'h002A;
        rom[9][74] = 16'h0009;
        rom[9][75] = 16'hFFDC;
        rom[9][76] = 16'h001D;
        rom[9][77] = 16'hFFC5;
        rom[9][78] = 16'hFFFC;
        rom[9][79] = 16'hFFF8;
        rom[9][80] = 16'h0037;
        rom[9][81] = 16'h000B;
        rom[9][82] = 16'h0042;
        rom[9][83] = 16'h000B;
        rom[9][84] = 16'h0007;
        rom[9][85] = 16'hFFC3;
        rom[9][86] = 16'hFFC6;
        rom[9][87] = 16'h0005;
        rom[9][88] = 16'hFFCF;
        rom[9][89] = 16'hFFF1;
        rom[9][90] = 16'h000E;
        rom[9][91] = 16'hFFC2;
        rom[9][92] = 16'h0015;
        rom[9][93] = 16'hFFDD;
        rom[9][94] = 16'hFFAB;
        rom[9][95] = 16'hFFE5;
        rom[9][96] = 16'hFFFF;
        rom[9][97] = 16'h000B;
        rom[9][98] = 16'hFFFC;
        rom[9][99] = 16'hFFEF;
        rom[9][100] = 16'hFFE2;
        rom[9][101] = 16'hFFFC;
        rom[9][102] = 16'h0034;
        rom[9][103] = 16'h001C;
        rom[9][104] = 16'hFFC6;
        rom[9][105] = 16'h0002;
        rom[9][106] = 16'hFFFE;
        rom[9][107] = 16'hFFF6;
        rom[9][108] = 16'hFFE9;
        rom[9][109] = 16'hFFFE;
        rom[9][110] = 16'h0039;
        rom[9][111] = 16'h0012;
        rom[9][112] = 16'hFFF2;
        rom[9][113] = 16'h0017;
        rom[9][114] = 16'h000A;
        rom[9][115] = 16'h0011;
        rom[9][116] = 16'hFFEC;
        rom[9][117] = 16'h001E;
        rom[9][118] = 16'hFFFE;
        rom[9][119] = 16'h0024;
        rom[9][120] = 16'hFFF0;
        rom[9][121] = 16'hFFB9;
        rom[9][122] = 16'h0012;
        rom[9][123] = 16'h0017;
        rom[9][124] = 16'hFFEA;
        rom[9][125] = 16'hFFEF;
        rom[9][126] = 16'hFFB7;
        rom[9][127] = 16'hFFD4;
        rom[10][0] = 16'hFFF7;
        rom[10][1] = 16'h0016;
        rom[10][2] = 16'hFFE6;
        rom[10][3] = 16'hFFBF;
        rom[10][4] = 16'h000C;
        rom[10][5] = 16'h001B;
        rom[10][6] = 16'h0019;
        rom[10][7] = 16'h0028;
        rom[10][8] = 16'h0012;
        rom[10][9] = 16'hFFC5;
        rom[10][10] = 16'h0024;
        rom[10][11] = 16'h0002;
        rom[10][12] = 16'hFFE5;
        rom[10][13] = 16'hFFDF;
        rom[10][14] = 16'h0016;
        rom[10][15] = 16'hFFC5;
        rom[10][16] = 16'h002E;
        rom[10][17] = 16'hFFED;
        rom[10][18] = 16'hFFFE;
        rom[10][19] = 16'h0013;
        rom[10][20] = 16'hFFE1;
        rom[10][21] = 16'hFFD2;
        rom[10][22] = 16'h001F;
        rom[10][23] = 16'hFFF6;
        rom[10][24] = 16'hFFCE;
        rom[10][25] = 16'h0017;
        rom[10][26] = 16'h001F;
        rom[10][27] = 16'h0023;
        rom[10][28] = 16'hFFFE;
        rom[10][29] = 16'hFFC9;
        rom[10][30] = 16'h0018;
        rom[10][31] = 16'hFFDB;
        rom[10][32] = 16'h0006;
        rom[10][33] = 16'h0010;
        rom[10][34] = 16'h0038;
        rom[10][35] = 16'hFFE9;
        rom[10][36] = 16'hFFEA;
        rom[10][37] = 16'hFFCB;
        rom[10][38] = 16'h0008;
        rom[10][39] = 16'hFFEF;
        rom[10][40] = 16'hFFD3;
        rom[10][41] = 16'hFFF7;
        rom[10][42] = 16'hFFDA;
        rom[10][43] = 16'hFFF5;
        rom[10][44] = 16'hFFE6;
        rom[10][45] = 16'hFFD7;
        rom[10][46] = 16'hFFF6;
        rom[10][47] = 16'hFFF7;
        rom[10][48] = 16'hFFE2;
        rom[10][49] = 16'h0038;
        rom[10][50] = 16'h0001;
        rom[10][51] = 16'hFFF5;
        rom[10][52] = 16'h0006;
        rom[10][53] = 16'hFFDF;
        rom[10][54] = 16'hFFCD;
        rom[10][55] = 16'hFFDD;
        rom[10][56] = 16'hFFF0;
        rom[10][57] = 16'hFFB8;
        rom[10][58] = 16'hFFDA;
        rom[10][59] = 16'h0007;
        rom[10][60] = 16'hFFF1;
        rom[10][61] = 16'hFFE6;
        rom[10][62] = 16'h0031;
        rom[10][63] = 16'hFFE9;
        rom[10][64] = 16'hFFDC;
        rom[10][65] = 16'hFFFB;
        rom[10][66] = 16'h0002;
        rom[10][67] = 16'h0029;
        rom[10][68] = 16'h0006;
        rom[10][69] = 16'h0009;
        rom[10][70] = 16'hFFD6;
        rom[10][71] = 16'h0024;
        rom[10][72] = 16'h0002;
        rom[10][73] = 16'hFFF3;
        rom[10][74] = 16'hFFC2;
        rom[10][75] = 16'hFFE6;
        rom[10][76] = 16'hFFCD;
        rom[10][77] = 16'hFFFE;
        rom[10][78] = 16'hFFEA;
        rom[10][79] = 16'hFFF4;
        rom[10][80] = 16'h0033;
        rom[10][81] = 16'hFFDB;
        rom[10][82] = 16'h001C;
        rom[10][83] = 16'hFFC4;
        rom[10][84] = 16'h0026;
        rom[10][85] = 16'h001A;
        rom[10][86] = 16'hFFF0;
        rom[10][87] = 16'h0022;
        rom[10][88] = 16'hFFE4;
        rom[10][89] = 16'hFFE1;
        rom[10][90] = 16'h0011;
        rom[10][91] = 16'h001E;
        rom[10][92] = 16'hFFFB;
        rom[10][93] = 16'hFFFA;
        rom[10][94] = 16'h0013;
        rom[10][95] = 16'hFFDE;
        rom[10][96] = 16'hFFF3;
        rom[10][97] = 16'h0013;
        rom[10][98] = 16'h0024;
        rom[10][99] = 16'hFFF9;
        rom[10][100] = 16'h0022;
        rom[10][101] = 16'hFFE6;
        rom[10][102] = 16'h001F;
        rom[10][103] = 16'hFFD9;
        rom[10][104] = 16'hFFE7;
        rom[10][105] = 16'h0029;
        rom[10][106] = 16'hFFCD;
        rom[10][107] = 16'h0015;
        rom[10][108] = 16'h001E;
        rom[10][109] = 16'hFFE7;
        rom[10][110] = 16'h000B;
        rom[10][111] = 16'hFFE3;
        rom[10][112] = 16'h002A;
        rom[10][113] = 16'hFFFB;
        rom[10][114] = 16'h0010;
        rom[10][115] = 16'hFFD3;
        rom[10][116] = 16'h0021;
        rom[10][117] = 16'h000C;
        rom[10][118] = 16'h001B;
        rom[10][119] = 16'hFFBE;
        rom[10][120] = 16'hFFFD;
        rom[10][121] = 16'h001F;
        rom[10][122] = 16'hFFFF;
        rom[10][123] = 16'h0021;
        rom[10][124] = 16'h0007;
        rom[10][125] = 16'hFFF1;
        rom[10][126] = 16'h0020;
        rom[10][127] = 16'h002A;
        rom[11][0] = 16'hFFE5;
        rom[11][1] = 16'h001F;
        rom[11][2] = 16'h0014;
        rom[11][3] = 16'hFFFD;
        rom[11][4] = 16'hFFEF;
        rom[11][5] = 16'h0018;
        rom[11][6] = 16'hFFEA;
        rom[11][7] = 16'h0019;
        rom[11][8] = 16'h0010;
        rom[11][9] = 16'h000F;
        rom[11][10] = 16'h000F;
        rom[11][11] = 16'hFFFA;
        rom[11][12] = 16'hFFBC;
        rom[11][13] = 16'hFFF4;
        rom[11][14] = 16'h002D;
        rom[11][15] = 16'h0012;
        rom[11][16] = 16'hFFED;
        rom[11][17] = 16'h0019;
        rom[11][18] = 16'hFFEF;
        rom[11][19] = 16'h0008;
        rom[11][20] = 16'h0008;
        rom[11][21] = 16'hFFFA;
        rom[11][22] = 16'h0019;
        rom[11][23] = 16'h000C;
        rom[11][24] = 16'h0015;
        rom[11][25] = 16'hFFFA;
        rom[11][26] = 16'h0025;
        rom[11][27] = 16'hFFFE;
        rom[11][28] = 16'hFFEC;
        rom[11][29] = 16'hFFFE;
        rom[11][30] = 16'hFFE6;
        rom[11][31] = 16'h0018;
        rom[11][32] = 16'hFFFF;
        rom[11][33] = 16'hFFEF;
        rom[11][34] = 16'hFFB5;
        rom[11][35] = 16'hFFE9;
        rom[11][36] = 16'h0024;
        rom[11][37] = 16'hFFDE;
        rom[11][38] = 16'h0016;
        rom[11][39] = 16'hFFFE;
        rom[11][40] = 16'h0007;
        rom[11][41] = 16'hFFFF;
        rom[11][42] = 16'h0029;
        rom[11][43] = 16'hFFB1;
        rom[11][44] = 16'hFFFA;
        rom[11][45] = 16'hFFF4;
        rom[11][46] = 16'h000A;
        rom[11][47] = 16'hFFC3;
        rom[11][48] = 16'hFFF5;
        rom[11][49] = 16'hFFE3;
        rom[11][50] = 16'h0011;
        rom[11][51] = 16'hFFD2;
        rom[11][52] = 16'hFFD2;
        rom[11][53] = 16'hFFF3;
        rom[11][54] = 16'hFFDA;
        rom[11][55] = 16'hFFEF;
        rom[11][56] = 16'hFFF3;
        rom[11][57] = 16'h0003;
        rom[11][58] = 16'hFFDC;
        rom[11][59] = 16'h0027;
        rom[11][60] = 16'hFFF3;
        rom[11][61] = 16'hFFF9;
        rom[11][62] = 16'h001B;
        rom[11][63] = 16'h000C;
        rom[11][64] = 16'hFFD7;
        rom[11][65] = 16'hFFEB;
        rom[11][66] = 16'h0001;
        rom[11][67] = 16'hFFE0;
        rom[11][68] = 16'hFFEF;
        rom[11][69] = 16'h0008;
        rom[11][70] = 16'h0027;
        rom[11][71] = 16'hFFA7;
        rom[11][72] = 16'hFFFD;
        rom[11][73] = 16'h0018;
        rom[11][74] = 16'h000C;
        rom[11][75] = 16'hFFFA;
        rom[11][76] = 16'hFFE1;
        rom[11][77] = 16'h0005;
        rom[11][78] = 16'h0016;
        rom[11][79] = 16'hFFCB;
        rom[11][80] = 16'h0046;
        rom[11][81] = 16'hFFE6;
        rom[11][82] = 16'h0014;
        rom[11][83] = 16'h001B;
        rom[11][84] = 16'h0016;
        rom[11][85] = 16'hFFEF;
        rom[11][86] = 16'h000C;
        rom[11][87] = 16'hFFC3;
        rom[11][88] = 16'hFFE4;
        rom[11][89] = 16'hFFEA;
        rom[11][90] = 16'hFFEC;
        rom[11][91] = 16'hFFE7;
        rom[11][92] = 16'h0004;
        rom[11][93] = 16'hFFDD;
        rom[11][94] = 16'hFFF8;
        rom[11][95] = 16'h0007;
        rom[11][96] = 16'hFFD0;
        rom[11][97] = 16'hFFB8;
        rom[11][98] = 16'hFFCC;
        rom[11][99] = 16'hFFF0;
        rom[11][100] = 16'h001F;
        rom[11][101] = 16'hFFF0;
        rom[11][102] = 16'hFFC9;
        rom[11][103] = 16'hFFE0;
        rom[11][104] = 16'hFFD6;
        rom[11][105] = 16'h002F;
        rom[11][106] = 16'h0005;
        rom[11][107] = 16'hFFE5;
        rom[11][108] = 16'h0008;
        rom[11][109] = 16'hFFCC;
        rom[11][110] = 16'hFFF3;
        rom[11][111] = 16'hFFFB;
        rom[11][112] = 16'hFFEA;
        rom[11][113] = 16'hFFE0;
        rom[11][114] = 16'hFFD2;
        rom[11][115] = 16'hFFB5;
        rom[11][116] = 16'hFFFE;
        rom[11][117] = 16'h0007;
        rom[11][118] = 16'h0012;
        rom[11][119] = 16'h0004;
        rom[11][120] = 16'hFFD5;
        rom[11][121] = 16'h0011;
        rom[11][122] = 16'hFFF4;
        rom[11][123] = 16'hFFF9;
        rom[11][124] = 16'hFFE8;
        rom[11][125] = 16'hFFC8;
        rom[11][126] = 16'hFFF0;
        rom[11][127] = 16'h000B;
        rom[12][0] = 16'h001C;
        rom[12][1] = 16'h0019;
        rom[12][2] = 16'h0039;
        rom[12][3] = 16'h0002;
        rom[12][4] = 16'hFFFE;
        rom[12][5] = 16'h0005;
        rom[12][6] = 16'h0004;
        rom[12][7] = 16'hFFE5;
        rom[12][8] = 16'hFFF4;
        rom[12][9] = 16'h0000;
        rom[12][10] = 16'hFFF7;
        rom[12][11] = 16'h0018;
        rom[12][12] = 16'h0038;
        rom[12][13] = 16'hFFF1;
        rom[12][14] = 16'hFFF4;
        rom[12][15] = 16'h0007;
        rom[12][16] = 16'h0021;
        rom[12][17] = 16'hFFD5;
        rom[12][18] = 16'h0039;
        rom[12][19] = 16'h0017;
        rom[12][20] = 16'h001E;
        rom[12][21] = 16'h0012;
        rom[12][22] = 16'hFFBC;
        rom[12][23] = 16'hFFDD;
        rom[12][24] = 16'hFFD8;
        rom[12][25] = 16'hFFF7;
        rom[12][26] = 16'h000A;
        rom[12][27] = 16'hFFDC;
        rom[12][28] = 16'hFFE4;
        rom[12][29] = 16'h0023;
        rom[12][30] = 16'hFFE5;
        rom[12][31] = 16'h0002;
        rom[12][32] = 16'h0042;
        rom[12][33] = 16'hFFE4;
        rom[12][34] = 16'hFFF4;
        rom[12][35] = 16'hFFC2;
        rom[12][36] = 16'h002F;
        rom[12][37] = 16'h0016;
        rom[12][38] = 16'hFFBF;
        rom[12][39] = 16'hFFDF;
        rom[12][40] = 16'h0006;
        rom[12][41] = 16'h0018;
        rom[12][42] = 16'hFFE1;
        rom[12][43] = 16'h000C;
        rom[12][44] = 16'h0004;
        rom[12][45] = 16'h0014;
        rom[12][46] = 16'hFFF8;
        rom[12][47] = 16'hFFFF;
        rom[12][48] = 16'hFFFC;
        rom[12][49] = 16'h0011;
        rom[12][50] = 16'hFFFA;
        rom[12][51] = 16'h0032;
        rom[12][52] = 16'h0015;
        rom[12][53] = 16'h001E;
        rom[12][54] = 16'hFFDD;
        rom[12][55] = 16'hFFEF;
        rom[12][56] = 16'h0029;
        rom[12][57] = 16'h0027;
        rom[12][58] = 16'h0002;
        rom[12][59] = 16'hFFF6;
        rom[12][60] = 16'hFFFE;
        rom[12][61] = 16'h002B;
        rom[12][62] = 16'h000A;
        rom[12][63] = 16'hFFF1;
        rom[12][64] = 16'h0030;
        rom[12][65] = 16'h0007;
        rom[12][66] = 16'h0012;
        rom[12][67] = 16'h0027;
        rom[12][68] = 16'h000E;
        rom[12][69] = 16'hFFFC;
        rom[12][70] = 16'hFFFB;
        rom[12][71] = 16'h0000;
        rom[12][72] = 16'h000A;
        rom[12][73] = 16'h002E;
        rom[12][74] = 16'hFFFE;
        rom[12][75] = 16'hFFDD;
        rom[12][76] = 16'hFFFE;
        rom[12][77] = 16'hFFE6;
        rom[12][78] = 16'h0012;
        rom[12][79] = 16'h0022;
        rom[12][80] = 16'hFFD6;
        rom[12][81] = 16'h0006;
        rom[12][82] = 16'hFFFD;
        rom[12][83] = 16'h0000;
        rom[12][84] = 16'h000C;
        rom[12][85] = 16'hFFC2;
        rom[12][86] = 16'h0020;
        rom[12][87] = 16'hFFD9;
        rom[12][88] = 16'h000A;
        rom[12][89] = 16'h0002;
        rom[12][90] = 16'h0023;
        rom[12][91] = 16'h0012;
        rom[12][92] = 16'hFFBA;
        rom[12][93] = 16'h0001;
        rom[12][94] = 16'h0016;
        rom[12][95] = 16'hFFE8;
        rom[12][96] = 16'hFFF7;
        rom[12][97] = 16'h0020;
        rom[12][98] = 16'h0027;
        rom[12][99] = 16'hFFF8;
        rom[12][100] = 16'hFFF4;
        rom[12][101] = 16'hFFF4;
        rom[12][102] = 16'h0010;
        rom[12][103] = 16'hFFFF;
        rom[12][104] = 16'h0016;
        rom[12][105] = 16'hFFE6;
        rom[12][106] = 16'h000C;
        rom[12][107] = 16'h0011;
        rom[12][108] = 16'h0022;
        rom[12][109] = 16'hFFD1;
        rom[12][110] = 16'hFFFE;
        rom[12][111] = 16'h0015;
        rom[12][112] = 16'hFFE5;
        rom[12][113] = 16'h003D;
        rom[12][114] = 16'h0032;
        rom[12][115] = 16'h0001;
        rom[12][116] = 16'hFFE2;
        rom[12][117] = 16'hFFF4;
        rom[12][118] = 16'hFFCA;
        rom[12][119] = 16'hFFFE;
        rom[12][120] = 16'hFFFD;
        rom[12][121] = 16'hFFEC;
        rom[12][122] = 16'hFFF9;
        rom[12][123] = 16'hFFC0;
        rom[12][124] = 16'hFFCC;
        rom[12][125] = 16'h0033;
        rom[12][126] = 16'hFFC8;
        rom[12][127] = 16'h0016;
        rom[13][0] = 16'hFFD3;
        rom[13][1] = 16'hFFF0;
        rom[13][2] = 16'hFFE7;
        rom[13][3] = 16'h0008;
        rom[13][4] = 16'hFFEA;
        rom[13][5] = 16'h0007;
        rom[13][6] = 16'h000F;
        rom[13][7] = 16'hFFF3;
        rom[13][8] = 16'hFFFF;
        rom[13][9] = 16'h0017;
        rom[13][10] = 16'h0024;
        rom[13][11] = 16'h0002;
        rom[13][12] = 16'h0017;
        rom[13][13] = 16'hFFD2;
        rom[13][14] = 16'h0002;
        rom[13][15] = 16'hFFCA;
        rom[13][16] = 16'hFFF0;
        rom[13][17] = 16'h0012;
        rom[13][18] = 16'hFFF6;
        rom[13][19] = 16'hFFF7;
        rom[13][20] = 16'h0010;
        rom[13][21] = 16'h0003;
        rom[13][22] = 16'hFFCA;
        rom[13][23] = 16'h0032;
        rom[13][24] = 16'hFFD4;
        rom[13][25] = 16'h0011;
        rom[13][26] = 16'h0016;
        rom[13][27] = 16'h001B;
        rom[13][28] = 16'h0007;
        rom[13][29] = 16'hFFDA;
        rom[13][30] = 16'h0017;
        rom[13][31] = 16'hFFD9;
        rom[13][32] = 16'h0007;
        rom[13][33] = 16'hFFEF;
        rom[13][34] = 16'h000B;
        rom[13][35] = 16'hFFD2;
        rom[13][36] = 16'hFFF2;
        rom[13][37] = 16'h0011;
        rom[13][38] = 16'hFFF5;
        rom[13][39] = 16'hFFEE;
        rom[13][40] = 16'hFFF5;
        rom[13][41] = 16'h0003;
        rom[13][42] = 16'h0010;
        rom[13][43] = 16'h0009;
        rom[13][44] = 16'h000A;
        rom[13][45] = 16'hFFF7;
        rom[13][46] = 16'h0016;
        rom[13][47] = 16'h0009;
        rom[13][48] = 16'hFFE4;
        rom[13][49] = 16'hFFF9;
        rom[13][50] = 16'h0007;
        rom[13][51] = 16'hFFD3;
        rom[13][52] = 16'hFFF4;
        rom[13][53] = 16'hFFEA;
        rom[13][54] = 16'hFFF6;
        rom[13][55] = 16'hFFE0;
        rom[13][56] = 16'hFFFC;
        rom[13][57] = 16'hFFC3;
        rom[13][58] = 16'h0003;
        rom[13][59] = 16'h0022;
        rom[13][60] = 16'hFFF8;
        rom[13][61] = 16'hFFFE;
        rom[13][62] = 16'h000C;
        rom[13][63] = 16'h0046;
        rom[13][64] = 16'hFFB2;
        rom[13][65] = 16'hFFB4;
        rom[13][66] = 16'h0013;
        rom[13][67] = 16'h0002;
        rom[13][68] = 16'hFFEB;
        rom[13][69] = 16'hFFD4;
        rom[13][70] = 16'hFFE2;
        rom[13][71] = 16'hFFF9;
        rom[13][72] = 16'hFFCD;
        rom[13][73] = 16'h0003;
        rom[13][74] = 16'hFFD9;
        rom[13][75] = 16'h0014;
        rom[13][76] = 16'h000C;
        rom[13][77] = 16'h001A;
        rom[13][78] = 16'hFFD2;
        rom[13][79] = 16'h0016;
        rom[13][80] = 16'h0018;
        rom[13][81] = 16'hFFE3;
        rom[13][82] = 16'h0020;
        rom[13][83] = 16'hFFFD;
        rom[13][84] = 16'hFFBF;
        rom[13][85] = 16'hFFFE;
        rom[13][86] = 16'hFFEF;
        rom[13][87] = 16'hFFFE;
        rom[13][88] = 16'h001D;
        rom[13][89] = 16'hFFF7;
        rom[13][90] = 16'h0032;
        rom[13][91] = 16'h0001;
        rom[13][92] = 16'hFFF4;
        rom[13][93] = 16'hFFDB;
        rom[13][94] = 16'hFFF5;
        rom[13][95] = 16'hFFBE;
        rom[13][96] = 16'hFFF0;
        rom[13][97] = 16'hFFF7;
        rom[13][98] = 16'h0029;
        rom[13][99] = 16'hFFDA;
        rom[13][100] = 16'h0024;
        rom[13][101] = 16'hFFCF;
        rom[13][102] = 16'h0001;
        rom[13][103] = 16'hFFE2;
        rom[13][104] = 16'h0005;
        rom[13][105] = 16'hFFB2;
        rom[13][106] = 16'hFFF8;
        rom[13][107] = 16'h000F;
        rom[13][108] = 16'hFFE0;
        rom[13][109] = 16'hFFC9;
        rom[13][110] = 16'hFFD5;
        rom[13][111] = 16'hFFBF;
        rom[13][112] = 16'hFFFC;
        rom[13][113] = 16'hFFF5;
        rom[13][114] = 16'hFFDE;
        rom[13][115] = 16'hFFD6;
        rom[13][116] = 16'h0014;
        rom[13][117] = 16'h0001;
        rom[13][118] = 16'h0024;
        rom[13][119] = 16'hFFDC;
        rom[13][120] = 16'h0004;
        rom[13][121] = 16'h000A;
        rom[13][122] = 16'h0029;
        rom[13][123] = 16'h0008;
        rom[13][124] = 16'hFFF5;
        rom[13][125] = 16'h003A;
        rom[13][126] = 16'h0019;
        rom[13][127] = 16'hFFF1;
        rom[14][0] = 16'h0013;
        rom[14][1] = 16'h0017;
        rom[14][2] = 16'hFFE5;
        rom[14][3] = 16'h0012;
        rom[14][4] = 16'h0011;
        rom[14][5] = 16'hFFE6;
        rom[14][6] = 16'hFFD6;
        rom[14][7] = 16'hFFD7;
        rom[14][8] = 16'h000C;
        rom[14][9] = 16'hFFE7;
        rom[14][10] = 16'h001D;
        rom[14][11] = 16'hFFE3;
        rom[14][12] = 16'hFFD4;
        rom[14][13] = 16'hFFDA;
        rom[14][14] = 16'hFFF7;
        rom[14][15] = 16'h000F;
        rom[14][16] = 16'hFFD2;
        rom[14][17] = 16'h001A;
        rom[14][18] = 16'h0011;
        rom[14][19] = 16'h0006;
        rom[14][20] = 16'h0013;
        rom[14][21] = 16'hFFFA;
        rom[14][22] = 16'hFFEA;
        rom[14][23] = 16'hFFD2;
        rom[14][24] = 16'hFFFE;
        rom[14][25] = 16'h0017;
        rom[14][26] = 16'h0032;
        rom[14][27] = 16'h0002;
        rom[14][28] = 16'hFFF9;
        rom[14][29] = 16'h0016;
        rom[14][30] = 16'hFFF9;
        rom[14][31] = 16'hFFC3;
        rom[14][32] = 16'hFFF9;
        rom[14][33] = 16'h000D;
        rom[14][34] = 16'hFFE3;
        rom[14][35] = 16'h0007;
        rom[14][36] = 16'hFFCB;
        rom[14][37] = 16'h0011;
        rom[14][38] = 16'h0015;
        rom[14][39] = 16'h0006;
        rom[14][40] = 16'hFFD4;
        rom[14][41] = 16'h0038;
        rom[14][42] = 16'h0003;
        rom[14][43] = 16'h001E;
        rom[14][44] = 16'hFFF4;
        rom[14][45] = 16'hFFF8;
        rom[14][46] = 16'hFFD2;
        rom[14][47] = 16'h000F;
        rom[14][48] = 16'hFFD9;
        rom[14][49] = 16'hFFE7;
        rom[14][50] = 16'h000C;
        rom[14][51] = 16'h0037;
        rom[14][52] = 16'hFFE9;
        rom[14][53] = 16'hFFBC;
        rom[14][54] = 16'h0010;
        rom[14][55] = 16'h000C;
        rom[14][56] = 16'h0010;
        rom[14][57] = 16'hFFC8;
        rom[14][58] = 16'hFFE3;
        rom[14][59] = 16'h0008;
        rom[14][60] = 16'hFFFD;
        rom[14][61] = 16'hFFF3;
        rom[14][62] = 16'hFFF6;
        rom[14][63] = 16'hFFFE;
        rom[14][64] = 16'h001B;
        rom[14][65] = 16'hFFF9;
        rom[14][66] = 16'hFFF2;
        rom[14][67] = 16'hFFF2;
        rom[14][68] = 16'hFFED;
        rom[14][69] = 16'hFFD0;
        rom[14][70] = 16'h0002;
        rom[14][71] = 16'hFFFD;
        rom[14][72] = 16'hFFB2;
        rom[14][73] = 16'h000B;
        rom[14][74] = 16'hFFCD;
        rom[14][75] = 16'hFFF9;
        rom[14][76] = 16'h001E;
        rom[14][77] = 16'hFFE7;
        rom[14][78] = 16'h001B;
        rom[14][79] = 16'hFFD8;
        rom[14][80] = 16'h000E;
        rom[14][81] = 16'hFFE8;
        rom[14][82] = 16'h001F;
        rom[14][83] = 16'h0002;
        rom[14][84] = 16'hFFBF;
        rom[14][85] = 16'hFFFD;
        rom[14][86] = 16'h001D;
        rom[14][87] = 16'hFFE0;
        rom[14][88] = 16'h0033;
        rom[14][89] = 16'h0026;
        rom[14][90] = 16'h0003;
        rom[14][91] = 16'hFFEA;
        rom[14][92] = 16'h0005;
        rom[14][93] = 16'h0003;
        rom[14][94] = 16'hFFC6;
        rom[14][95] = 16'h0021;
        rom[14][96] = 16'h000A;
        rom[14][97] = 16'h0002;
        rom[14][98] = 16'hFFF6;
        rom[14][99] = 16'hFFF4;
        rom[14][100] = 16'hFFE7;
        rom[14][101] = 16'h0014;
        rom[14][102] = 16'hFFEC;
        rom[14][103] = 16'hFFD6;
        rom[14][104] = 16'h0016;
        rom[14][105] = 16'hFFE7;
        rom[14][106] = 16'hFFFE;
        rom[14][107] = 16'hFFEA;
        rom[14][108] = 16'hFFD4;
        rom[14][109] = 16'h0002;
        rom[14][110] = 16'hFFFA;
        rom[14][111] = 16'hFFF4;
        rom[14][112] = 16'hFFDF;
        rom[14][113] = 16'h0012;
        rom[14][114] = 16'hFFF5;
        rom[14][115] = 16'hFFE3;
        rom[14][116] = 16'hFFF5;
        rom[14][117] = 16'hFFFE;
        rom[14][118] = 16'hFFF5;
        rom[14][119] = 16'hFFFB;
        rom[14][120] = 16'hFFE0;
        rom[14][121] = 16'hFFF2;
        rom[14][122] = 16'hFFB7;
        rom[14][123] = 16'h0007;
        rom[14][124] = 16'hFFC9;
        rom[14][125] = 16'h0005;
        rom[14][126] = 16'hFFE5;
        rom[14][127] = 16'hFFCD;
        rom[15][0] = 16'hFFFD;
        rom[15][1] = 16'h0029;
        rom[15][2] = 16'hFFFC;
        rom[15][3] = 16'h000B;
        rom[15][4] = 16'hFFF6;
        rom[15][5] = 16'h001A;
        rom[15][6] = 16'h001A;
        rom[15][7] = 16'hFFEE;
        rom[15][8] = 16'h0006;
        rom[15][9] = 16'hFFEF;
        rom[15][10] = 16'hFFFD;
        rom[15][11] = 16'h000A;
        rom[15][12] = 16'hFFC3;
        rom[15][13] = 16'hFFE7;
        rom[15][14] = 16'hFFEE;
        rom[15][15] = 16'hFFEF;
        rom[15][16] = 16'h0001;
        rom[15][17] = 16'hFFD9;
        rom[15][18] = 16'hFFF4;
        rom[15][19] = 16'h0016;
        rom[15][20] = 16'hFFFD;
        rom[15][21] = 16'h0019;
        rom[15][22] = 16'hFFF4;
        rom[15][23] = 16'h0029;
        rom[15][24] = 16'h0006;
        rom[15][25] = 16'h0023;
        rom[15][26] = 16'hFFD6;
        rom[15][27] = 16'hFFE5;
        rom[15][28] = 16'hFFEE;
        rom[15][29] = 16'hFFD7;
        rom[15][30] = 16'h0011;
        rom[15][31] = 16'hFFE3;
        rom[15][32] = 16'hFFFC;
        rom[15][33] = 16'hFFDE;
        rom[15][34] = 16'h000F;
        rom[15][35] = 16'hFFB7;
        rom[15][36] = 16'hFFE5;
        rom[15][37] = 16'h0002;
        rom[15][38] = 16'hFFFE;
        rom[15][39] = 16'hFFE2;
        rom[15][40] = 16'hFFBF;
        rom[15][41] = 16'h0015;
        rom[15][42] = 16'hFFEA;
        rom[15][43] = 16'hFFC2;
        rom[15][44] = 16'hFFF8;
        rom[15][45] = 16'hFFE1;
        rom[15][46] = 16'h0012;
        rom[15][47] = 16'hFFD4;
        rom[15][48] = 16'hFFCF;
        rom[15][49] = 16'hFFD1;
        rom[15][50] = 16'h0019;
        rom[15][51] = 16'hFFF6;
        rom[15][52] = 16'h000B;
        rom[15][53] = 16'hFFBC;
        rom[15][54] = 16'hFFF4;
        rom[15][55] = 16'hFFFB;
        rom[15][56] = 16'hFFD2;
        rom[15][57] = 16'hFFD5;
        rom[15][58] = 16'h0016;
        rom[15][59] = 16'h0027;
        rom[15][60] = 16'hFFF5;
        rom[15][61] = 16'hFFEE;
        rom[15][62] = 16'hFFFE;
        rom[15][63] = 16'h0009;
        rom[15][64] = 16'hFFE5;
        rom[15][65] = 16'hFFF6;
        rom[15][66] = 16'h0007;
        rom[15][67] = 16'hFFEE;
        rom[15][68] = 16'hFFCE;
        rom[15][69] = 16'h000E;
        rom[15][70] = 16'h000D;
        rom[15][71] = 16'h0002;
        rom[15][72] = 16'h000A;
        rom[15][73] = 16'hFFD5;
        rom[15][74] = 16'hFFD5;
        rom[15][75] = 16'h0021;
        rom[15][76] = 16'h000C;
        rom[15][77] = 16'hFFFE;
        rom[15][78] = 16'h0006;
        rom[15][79] = 16'hFFF9;
        rom[15][80] = 16'h0011;
        rom[15][81] = 16'h000C;
        rom[15][82] = 16'h003D;
        rom[15][83] = 16'hFFE0;
        rom[15][84] = 16'hFFC8;
        rom[15][85] = 16'h0007;
        rom[15][86] = 16'hFFF4;
        rom[15][87] = 16'h0009;
        rom[15][88] = 16'h0004;
        rom[15][89] = 16'hFFFE;
        rom[15][90] = 16'h0025;
        rom[15][91] = 16'h001F;
        rom[15][92] = 16'h002B;
        rom[15][93] = 16'h000E;
        rom[15][94] = 16'h0009;
        rom[15][95] = 16'hFFD9;
        rom[15][96] = 16'h0000;
        rom[15][97] = 16'h0018;
        rom[15][98] = 16'h0024;
        rom[15][99] = 16'hFFE5;
        rom[15][100] = 16'h0021;
        rom[15][101] = 16'h0038;
        rom[15][102] = 16'hFFDB;
        rom[15][103] = 16'hFFE1;
        rom[15][104] = 16'h0007;
        rom[15][105] = 16'h0004;
        rom[15][106] = 16'hFFFF;
        rom[15][107] = 16'hFFF9;
        rom[15][108] = 16'hFFFE;
        rom[15][109] = 16'hFF98;
        rom[15][110] = 16'h0021;
        rom[15][111] = 16'h001A;
        rom[15][112] = 16'hFFDF;
        rom[15][113] = 16'h0002;
        rom[15][114] = 16'hFFE0;
        rom[15][115] = 16'hFFF2;
        rom[15][116] = 16'h000D;
        rom[15][117] = 16'h0036;
        rom[15][118] = 16'h0026;
        rom[15][119] = 16'h0003;
        rom[15][120] = 16'h0006;
        rom[15][121] = 16'h0016;
        rom[15][122] = 16'h001D;
        rom[15][123] = 16'h0000;
        rom[15][124] = 16'h000A;
        rom[15][125] = 16'h0022;
        rom[15][126] = 16'hFFE3;
        rom[15][127] = 16'h0029;
        rom[16][0] = 16'hFFFA;
        rom[16][1] = 16'h001D;
        rom[16][2] = 16'hFFC0;
        rom[16][3] = 16'h0027;
        rom[16][4] = 16'h0002;
        rom[16][5] = 16'hFFDE;
        rom[16][6] = 16'h0017;
        rom[16][7] = 16'hFFD7;
        rom[16][8] = 16'h000C;
        rom[16][9] = 16'hFFD7;
        rom[16][10] = 16'h0016;
        rom[16][11] = 16'hFFE7;
        rom[16][12] = 16'h0012;
        rom[16][13] = 16'hFFE3;
        rom[16][14] = 16'h000C;
        rom[16][15] = 16'h0015;
        rom[16][16] = 16'h000E;
        rom[16][17] = 16'hFFD1;
        rom[16][18] = 16'hFFEB;
        rom[16][19] = 16'h001B;
        rom[16][20] = 16'h0014;
        rom[16][21] = 16'h0029;
        rom[16][22] = 16'hFFE2;
        rom[16][23] = 16'h000B;
        rom[16][24] = 16'hFFFB;
        rom[16][25] = 16'hFFFC;
        rom[16][26] = 16'hFFF6;
        rom[16][27] = 16'h0008;
        rom[16][28] = 16'hFFFB;
        rom[16][29] = 16'h0022;
        rom[16][30] = 16'h0016;
        rom[16][31] = 16'h002D;
        rom[16][32] = 16'hFFA4;
        rom[16][33] = 16'h0003;
        rom[16][34] = 16'h000D;
        rom[16][35] = 16'hFFF9;
        rom[16][36] = 16'h002D;
        rom[16][37] = 16'h001A;
        rom[16][38] = 16'hFFCC;
        rom[16][39] = 16'h0024;
        rom[16][40] = 16'hFFFD;
        rom[16][41] = 16'hFFE8;
        rom[16][42] = 16'h0009;
        rom[16][43] = 16'hFFC3;
        rom[16][44] = 16'h0011;
        rom[16][45] = 16'hFFD5;
        rom[16][46] = 16'hFFF7;
        rom[16][47] = 16'h0011;
        rom[16][48] = 16'hFFFC;
        rom[16][49] = 16'hFFFE;
        rom[16][50] = 16'hFFD9;
        rom[16][51] = 16'hFFFA;
        rom[16][52] = 16'hFF96;
        rom[16][53] = 16'hFFDC;
        rom[16][54] = 16'h002E;
        rom[16][55] = 16'h0029;
        rom[16][56] = 16'hFFD2;
        rom[16][57] = 16'hFFE4;
        rom[16][58] = 16'h0017;
        rom[16][59] = 16'hFFF9;
        rom[16][60] = 16'h0020;
        rom[16][61] = 16'h0009;
        rom[16][62] = 16'h0007;
        rom[16][63] = 16'hFFF4;
        rom[16][64] = 16'h001D;
        rom[16][65] = 16'h0004;
        rom[16][66] = 16'hFFDB;
        rom[16][67] = 16'h0000;
        rom[16][68] = 16'hFFE3;
        rom[16][69] = 16'h001B;
        rom[16][70] = 16'hFFD3;
        rom[16][71] = 16'hFFBB;
        rom[16][72] = 16'h0014;
        rom[16][73] = 16'hFFFC;
        rom[16][74] = 16'h0007;
        rom[16][75] = 16'hFFF4;
        rom[16][76] = 16'h0014;
        rom[16][77] = 16'h0025;
        rom[16][78] = 16'h002E;
        rom[16][79] = 16'h0006;
        rom[16][80] = 16'hFFDA;
        rom[16][81] = 16'h000D;
        rom[16][82] = 16'hFFFC;
        rom[16][83] = 16'hFFF8;
        rom[16][84] = 16'hFFF5;
        rom[16][85] = 16'hFFEA;
        rom[16][86] = 16'h000F;
        rom[16][87] = 16'h0008;
        rom[16][88] = 16'hFFDC;
        rom[16][89] = 16'h002C;
        rom[16][90] = 16'hFFF5;
        rom[16][91] = 16'hFFEE;
        rom[16][92] = 16'h0024;
        rom[16][93] = 16'h000A;
        rom[16][94] = 16'hFFEC;
        rom[16][95] = 16'hFFEC;
        rom[16][96] = 16'hFFF4;
        rom[16][97] = 16'h0012;
        rom[16][98] = 16'h0023;
        rom[16][99] = 16'h000D;
        rom[16][100] = 16'h000E;
        rom[16][101] = 16'hFFE3;
        rom[16][102] = 16'hFFFB;
        rom[16][103] = 16'hFFDC;
        rom[16][104] = 16'hFFF3;
        rom[16][105] = 16'hFFF9;
        rom[16][106] = 16'hFFE2;
        rom[16][107] = 16'hFFC1;
        rom[16][108] = 16'hFFEE;
        rom[16][109] = 16'hFFFB;
        rom[16][110] = 16'h0007;
        rom[16][111] = 16'h0015;
        rom[16][112] = 16'hFFF3;
        rom[16][113] = 16'hFFF3;
        rom[16][114] = 16'hFFF4;
        rom[16][115] = 16'h001D;
        rom[16][116] = 16'h001B;
        rom[16][117] = 16'hFFFC;
        rom[16][118] = 16'hFFD4;
        rom[16][119] = 16'hFFD2;
        rom[16][120] = 16'h0002;
        rom[16][121] = 16'h000C;
        rom[16][122] = 16'h0003;
        rom[16][123] = 16'h0011;
        rom[16][124] = 16'h000F;
        rom[16][125] = 16'hFFFA;
        rom[16][126] = 16'hFFC3;
        rom[16][127] = 16'hFFDE;
        rom[17][0] = 16'hFFEF;
        rom[17][1] = 16'h0000;
        rom[17][2] = 16'hFFF6;
        rom[17][3] = 16'h0008;
        rom[17][4] = 16'h000F;
        rom[17][5] = 16'h001C;
        rom[17][6] = 16'h002E;
        rom[17][7] = 16'hFFEF;
        rom[17][8] = 16'hFFD8;
        rom[17][9] = 16'hFFA6;
        rom[17][10] = 16'hFFC9;
        rom[17][11] = 16'hFFD5;
        rom[17][12] = 16'hFFB1;
        rom[17][13] = 16'hFFC3;
        rom[17][14] = 16'h0004;
        rom[17][15] = 16'hFFF6;
        rom[17][16] = 16'h0007;
        rom[17][17] = 16'hFFCB;
        rom[17][18] = 16'hFFF9;
        rom[17][19] = 16'hFFEE;
        rom[17][20] = 16'hFFEA;
        rom[17][21] = 16'h0011;
        rom[17][22] = 16'h000D;
        rom[17][23] = 16'hFFFC;
        rom[17][24] = 16'hFFCE;
        rom[17][25] = 16'hFFE1;
        rom[17][26] = 16'h001F;
        rom[17][27] = 16'hFFDD;
        rom[17][28] = 16'hFFF4;
        rom[17][29] = 16'hFFC1;
        rom[17][30] = 16'hFFE2;
        rom[17][31] = 16'hFFDE;
        rom[17][32] = 16'hFFEC;
        rom[17][33] = 16'h0006;
        rom[17][34] = 16'hFFF9;
        rom[17][35] = 16'h0007;
        rom[17][36] = 16'h0015;
        rom[17][37] = 16'hFFE8;
        rom[17][38] = 16'hFFDC;
        rom[17][39] = 16'h0033;
        rom[17][40] = 16'hFFF5;
        rom[17][41] = 16'h0011;
        rom[17][42] = 16'h005A;
        rom[17][43] = 16'h0014;
        rom[17][44] = 16'h0015;
        rom[17][45] = 16'h0007;
        rom[17][46] = 16'h000C;
        rom[17][47] = 16'hFFCD;
        rom[17][48] = 16'h0009;
        rom[17][49] = 16'h0004;
        rom[17][50] = 16'h001B;
        rom[17][51] = 16'hFFD1;
        rom[17][52] = 16'h0019;
        rom[17][53] = 16'h0010;
        rom[17][54] = 16'h000A;
        rom[17][55] = 16'hFFFF;
        rom[17][56] = 16'hFFDF;
        rom[17][57] = 16'h002E;
        rom[17][58] = 16'hFFFE;
        rom[17][59] = 16'hFFB1;
        rom[17][60] = 16'h0024;
        rom[17][61] = 16'hFFD2;
        rom[17][62] = 16'h0003;
        rom[17][63] = 16'h002B;
        rom[17][64] = 16'hFFD0;
        rom[17][65] = 16'hFFFA;
        rom[17][66] = 16'hFFEC;
        rom[17][67] = 16'hFFF9;
        rom[17][68] = 16'h0033;
        rom[17][69] = 16'h0000;
        rom[17][70] = 16'hFFFF;
        rom[17][71] = 16'h002D;
        rom[17][72] = 16'hFFD0;
        rom[17][73] = 16'hFFEA;
        rom[17][74] = 16'h001D;
        rom[17][75] = 16'h0017;
        rom[17][76] = 16'hFFBA;
        rom[17][77] = 16'h0005;
        rom[17][78] = 16'h000B;
        rom[17][79] = 16'hFFE6;
        rom[17][80] = 16'hFFFC;
        rom[17][81] = 16'h0034;
        rom[17][82] = 16'h0024;
        rom[17][83] = 16'hFFD1;
        rom[17][84] = 16'h0037;
        rom[17][85] = 16'h002F;
        rom[17][86] = 16'hFFF3;
        rom[17][87] = 16'h0007;
        rom[17][88] = 16'h0004;
        rom[17][89] = 16'h001D;
        rom[17][90] = 16'hFFFE;
        rom[17][91] = 16'h000C;
        rom[17][92] = 16'hFFB8;
        rom[17][93] = 16'h001C;
        rom[17][94] = 16'hFFEE;
        rom[17][95] = 16'h0009;
        rom[17][96] = 16'h0019;
        rom[17][97] = 16'h001C;
        rom[17][98] = 16'hFFE1;
        rom[17][99] = 16'h002C;
        rom[17][100] = 16'hFFE7;
        rom[17][101] = 16'h001B;
        rom[17][102] = 16'h0032;
        rom[17][103] = 16'hFFE2;
        rom[17][104] = 16'h000F;
        rom[17][105] = 16'hFFF9;
        rom[17][106] = 16'hFFF6;
        rom[17][107] = 16'hFFF5;
        rom[17][108] = 16'hFFE4;
        rom[17][109] = 16'h0009;
        rom[17][110] = 16'hFFFA;
        rom[17][111] = 16'h001F;
        rom[17][112] = 16'hFFEE;
        rom[17][113] = 16'h0007;
        rom[17][114] = 16'h0016;
        rom[17][115] = 16'h002E;
        rom[17][116] = 16'h0006;
        rom[17][117] = 16'h000C;
        rom[17][118] = 16'h0017;
        rom[17][119] = 16'h0027;
        rom[17][120] = 16'hFFEA;
        rom[17][121] = 16'hFFF0;
        rom[17][122] = 16'hFFCE;
        rom[17][123] = 16'hFFD7;
        rom[17][124] = 16'h0020;
        rom[17][125] = 16'hFFF8;
        rom[17][126] = 16'hFFFA;
        rom[17][127] = 16'h0015;
        rom[18][0] = 16'h000F;
        rom[18][1] = 16'h0000;
        rom[18][2] = 16'hFFFB;
        rom[18][3] = 16'h002D;
        rom[18][4] = 16'h0012;
        rom[18][5] = 16'hFFDC;
        rom[18][6] = 16'h0011;
        rom[18][7] = 16'hFFEE;
        rom[18][8] = 16'hFFE1;
        rom[18][9] = 16'hFFCB;
        rom[18][10] = 16'hFFCD;
        rom[18][11] = 16'h0041;
        rom[18][12] = 16'hFFB9;
        rom[18][13] = 16'hFFE0;
        rom[18][14] = 16'hFFFD;
        rom[18][15] = 16'hFFB3;
        rom[18][16] = 16'h004B;
        rom[18][17] = 16'hFFF3;
        rom[18][18] = 16'h001B;
        rom[18][19] = 16'hFFE8;
        rom[18][20] = 16'h0027;
        rom[18][21] = 16'hFFD6;
        rom[18][22] = 16'hFFE3;
        rom[18][23] = 16'hFFFD;
        rom[18][24] = 16'h000E;
        rom[18][25] = 16'hFFEE;
        rom[18][26] = 16'h0011;
        rom[18][27] = 16'hFFFE;
        rom[18][28] = 16'hFFF5;
        rom[18][29] = 16'hFFD3;
        rom[18][30] = 16'hFFD2;
        rom[18][31] = 16'hFFE5;
        rom[18][32] = 16'h001C;
        rom[18][33] = 16'hFFD2;
        rom[18][34] = 16'hFFBF;
        rom[18][35] = 16'hFFF3;
        rom[18][36] = 16'h0010;
        rom[18][37] = 16'hFFEC;
        rom[18][38] = 16'hFFAA;
        rom[18][39] = 16'hFFE3;
        rom[18][40] = 16'hFFF1;
        rom[18][41] = 16'hFFF9;
        rom[18][42] = 16'hFFD1;
        rom[18][43] = 16'hFFF3;
        rom[18][44] = 16'hFFBB;
        rom[18][45] = 16'hFFEA;
        rom[18][46] = 16'h0036;
        rom[18][47] = 16'hFFCD;
        rom[18][48] = 16'h0012;
        rom[18][49] = 16'hFFFE;
        rom[18][50] = 16'h001B;
        rom[18][51] = 16'h001F;
        rom[18][52] = 16'hFFFB;
        rom[18][53] = 16'h0016;
        rom[18][54] = 16'h0024;
        rom[18][55] = 16'hFFB5;
        rom[18][56] = 16'hFFC4;
        rom[18][57] = 16'h004F;
        rom[18][58] = 16'hFFEE;
        rom[18][59] = 16'h0011;
        rom[18][60] = 16'h0001;
        rom[18][61] = 16'hFFC9;
        rom[18][62] = 16'hFFDB;
        rom[18][63] = 16'h0041;
        rom[18][64] = 16'hFFFF;
        rom[18][65] = 16'hFFEC;
        rom[18][66] = 16'hFFFA;
        rom[18][67] = 16'hFFF6;
        rom[18][68] = 16'hFFEB;
        rom[18][69] = 16'hFFCD;
        rom[18][70] = 16'hFFE5;
        rom[18][71] = 16'h001F;
        rom[18][72] = 16'h0031;
        rom[18][73] = 16'hFFC4;
        rom[18][74] = 16'h001F;
        rom[18][75] = 16'hFFE2;
        rom[18][76] = 16'h0006;
        rom[18][77] = 16'hFFD7;
        rom[18][78] = 16'hFFEE;
        rom[18][79] = 16'h0010;
        rom[18][80] = 16'hFFFD;
        rom[18][81] = 16'h0007;
        rom[18][82] = 16'h0033;
        rom[18][83] = 16'hFFA3;
        rom[18][84] = 16'hFFB5;
        rom[18][85] = 16'h0038;
        rom[18][86] = 16'h0007;
        rom[18][87] = 16'h0035;
        rom[18][88] = 16'hFFEE;
        rom[18][89] = 16'hFFF2;
        rom[18][90] = 16'h002E;
        rom[18][91] = 16'h0036;
        rom[18][92] = 16'h0000;
        rom[18][93] = 16'hFFDC;
        rom[18][94] = 16'hFFE5;
        rom[18][95] = 16'h0009;
        rom[18][96] = 16'h0010;
        rom[18][97] = 16'h0019;
        rom[18][98] = 16'hFFF0;
        rom[18][99] = 16'hFFEB;
        rom[18][100] = 16'hFFCB;
        rom[18][101] = 16'h0027;
        rom[18][102] = 16'h000B;
        rom[18][103] = 16'hFFFD;
        rom[18][104] = 16'hFFFE;
        rom[18][105] = 16'h0009;
        rom[18][106] = 16'hFFEF;
        rom[18][107] = 16'hFFC7;
        rom[18][108] = 16'h0000;
        rom[18][109] = 16'h0026;
        rom[18][110] = 16'hFFE4;
        rom[18][111] = 16'hFFF2;
        rom[18][112] = 16'h0014;
        rom[18][113] = 16'hFFEF;
        rom[18][114] = 16'h0023;
        rom[18][115] = 16'hFFFB;
        rom[18][116] = 16'hFFEE;
        rom[18][117] = 16'hFFE1;
        rom[18][118] = 16'hFFF4;
        rom[18][119] = 16'hFFEF;
        rom[18][120] = 16'h0002;
        rom[18][121] = 16'h000F;
        rom[18][122] = 16'h0026;
        rom[18][123] = 16'hFFCE;
        rom[18][124] = 16'h0023;
        rom[18][125] = 16'h0011;
        rom[18][126] = 16'hFFFB;
        rom[18][127] = 16'hFFF0;
        rom[19][0] = 16'hFFF3;
        rom[19][1] = 16'h0019;
        rom[19][2] = 16'h000C;
        rom[19][3] = 16'h0034;
        rom[19][4] = 16'hFFDC;
        rom[19][5] = 16'hFFF9;
        rom[19][6] = 16'hFFDA;
        rom[19][7] = 16'hFFF4;
        rom[19][8] = 16'hFFE7;
        rom[19][9] = 16'h002A;
        rom[19][10] = 16'h0001;
        rom[19][11] = 16'h0007;
        rom[19][12] = 16'hFFF1;
        rom[19][13] = 16'hFFC4;
        rom[19][14] = 16'h0007;
        rom[19][15] = 16'hFFFF;
        rom[19][16] = 16'hFFF3;
        rom[19][17] = 16'hFFE1;
        rom[19][18] = 16'hFFFD;
        rom[19][19] = 16'h0021;
        rom[19][20] = 16'h0011;
        rom[19][21] = 16'hFFFE;
        rom[19][22] = 16'h0008;
        rom[19][23] = 16'h001F;
        rom[19][24] = 16'hFFFE;
        rom[19][25] = 16'hFFEA;
        rom[19][26] = 16'h0002;
        rom[19][27] = 16'hFFE0;
        rom[19][28] = 16'h000F;
        rom[19][29] = 16'h0008;
        rom[19][30] = 16'hFFE6;
        rom[19][31] = 16'hFFCF;
        rom[19][32] = 16'h0025;
        rom[19][33] = 16'h0009;
        rom[19][34] = 16'hFF99;
        rom[19][35] = 16'h001E;
        rom[19][36] = 16'h000F;
        rom[19][37] = 16'h0007;
        rom[19][38] = 16'h0017;
        rom[19][39] = 16'h0015;
        rom[19][40] = 16'hFFEF;
        rom[19][41] = 16'h0012;
        rom[19][42] = 16'hFFF8;
        rom[19][43] = 16'h000A;
        rom[19][44] = 16'hFFF9;
        rom[19][45] = 16'h001B;
        rom[19][46] = 16'h002E;
        rom[19][47] = 16'hFFBB;
        rom[19][48] = 16'hFFDC;
        rom[19][49] = 16'hFFE6;
        rom[19][50] = 16'hFFF2;
        rom[19][51] = 16'hFFEE;
        rom[19][52] = 16'hFFFC;
        rom[19][53] = 16'h0019;
        rom[19][54] = 16'h001A;
        rom[19][55] = 16'hFFE6;
        rom[19][56] = 16'hFFE5;
        rom[19][57] = 16'hFFFF;
        rom[19][58] = 16'hFFD7;
        rom[19][59] = 16'hFFFF;
        rom[19][60] = 16'hFFF4;
        rom[19][61] = 16'hFFFB;
        rom[19][62] = 16'h001F;
        rom[19][63] = 16'hFFF0;
        rom[19][64] = 16'hFFFE;
        rom[19][65] = 16'hFFE1;
        rom[19][66] = 16'hFFEF;
        rom[19][67] = 16'hFFDC;
        rom[19][68] = 16'hFFE7;
        rom[19][69] = 16'hFFFC;
        rom[19][70] = 16'h0029;
        rom[19][71] = 16'h0007;
        rom[19][72] = 16'hFFFA;
        rom[19][73] = 16'hFFE0;
        rom[19][74] = 16'hFFDF;
        rom[19][75] = 16'h0011;
        rom[19][76] = 16'h0004;
        rom[19][77] = 16'hFFE1;
        rom[19][78] = 16'hFFF4;
        rom[19][79] = 16'h0016;
        rom[19][80] = 16'hFFE9;
        rom[19][81] = 16'h0022;
        rom[19][82] = 16'h0012;
        rom[19][83] = 16'h0010;
        rom[19][84] = 16'h000C;
        rom[19][85] = 16'hFFF3;
        rom[19][86] = 16'h001B;
        rom[19][87] = 16'hFFE5;
        rom[19][88] = 16'hFFE3;
        rom[19][89] = 16'h0013;
        rom[19][90] = 16'hFFF0;
        rom[19][91] = 16'h001B;
        rom[19][92] = 16'hFFB7;
        rom[19][93] = 16'h0022;
        rom[19][94] = 16'hFFC1;
        rom[19][95] = 16'h0001;
        rom[19][96] = 16'h000D;
        rom[19][97] = 16'hFFE9;
        rom[19][98] = 16'h001A;
        rom[19][99] = 16'hFFEC;
        rom[19][100] = 16'h002C;
        rom[19][101] = 16'h0029;
        rom[19][102] = 16'hFFE3;
        rom[19][103] = 16'h000B;
        rom[19][104] = 16'h0006;
        rom[19][105] = 16'hFFCE;
        rom[19][106] = 16'h000B;
        rom[19][107] = 16'h003A;
        rom[19][108] = 16'hFFEE;
        rom[19][109] = 16'h001A;
        rom[19][110] = 16'hFFE9;
        rom[19][111] = 16'h001C;
        rom[19][112] = 16'h000C;
        rom[19][113] = 16'h0010;
        rom[19][114] = 16'hFFF4;
        rom[19][115] = 16'hFFE2;
        rom[19][116] = 16'h0029;
        rom[19][117] = 16'h0024;
        rom[19][118] = 16'hFFE6;
        rom[19][119] = 16'h002D;
        rom[19][120] = 16'hFFFE;
        rom[19][121] = 16'h0018;
        rom[19][122] = 16'hFFFD;
        rom[19][123] = 16'h0063;
        rom[19][124] = 16'h0037;
        rom[19][125] = 16'hFFFC;
        rom[19][126] = 16'h0009;
        rom[19][127] = 16'h0002;
        rom[20][0] = 16'h0028;
        rom[20][1] = 16'hFFCB;
        rom[20][2] = 16'hFFAF;
        rom[20][3] = 16'hFFD0;
        rom[20][4] = 16'hFFFE;
        rom[20][5] = 16'h000F;
        rom[20][6] = 16'hFFD7;
        rom[20][7] = 16'h0022;
        rom[20][8] = 16'h001D;
        rom[20][9] = 16'hFFDC;
        rom[20][10] = 16'hFFED;
        rom[20][11] = 16'hFFBF;
        rom[20][12] = 16'h0008;
        rom[20][13] = 16'h002B;
        rom[20][14] = 16'h0015;
        rom[20][15] = 16'hFFE0;
        rom[20][16] = 16'hFFED;
        rom[20][17] = 16'h002B;
        rom[20][18] = 16'hFFEE;
        rom[20][19] = 16'hFFE5;
        rom[20][20] = 16'hFFEA;
        rom[20][21] = 16'hFFDC;
        rom[20][22] = 16'hFFF2;
        rom[20][23] = 16'h0030;
        rom[20][24] = 16'hFFFE;
        rom[20][25] = 16'hFFBF;
        rom[20][26] = 16'h0007;
        rom[20][27] = 16'hFFAC;
        rom[20][28] = 16'hFFF8;
        rom[20][29] = 16'h001F;
        rom[20][30] = 16'hFFFF;
        rom[20][31] = 16'h0019;
        rom[20][32] = 16'hFFD8;
        rom[20][33] = 16'h000C;
        rom[20][34] = 16'h0028;
        rom[20][35] = 16'hFFFF;
        rom[20][36] = 16'hFFC9;
        rom[20][37] = 16'hFFCE;
        rom[20][38] = 16'hFFDA;
        rom[20][39] = 16'h0002;
        rom[20][40] = 16'h001B;
        rom[20][41] = 16'hFFE4;
        rom[20][42] = 16'h000C;
        rom[20][43] = 16'h0012;
        rom[20][44] = 16'h001D;
        rom[20][45] = 16'hFFF1;
        rom[20][46] = 16'hFFE4;
        rom[20][47] = 16'h0004;
        rom[20][48] = 16'hFFEB;
        rom[20][49] = 16'h0025;
        rom[20][50] = 16'h0005;
        rom[20][51] = 16'h0057;
        rom[20][52] = 16'hFFE8;
        rom[20][53] = 16'h001A;
        rom[20][54] = 16'hFFD3;
        rom[20][55] = 16'hFFEF;
        rom[20][56] = 16'h0001;
        rom[20][57] = 16'h0027;
        rom[20][58] = 16'h0032;
        rom[20][59] = 16'hFFDD;
        rom[20][60] = 16'hFFFA;
        rom[20][61] = 16'h0062;
        rom[20][62] = 16'hFFCE;
        rom[20][63] = 16'h0014;
        rom[20][64] = 16'hFFEE;
        rom[20][65] = 16'h001B;
        rom[20][66] = 16'h0013;
        rom[20][67] = 16'hFFE1;
        rom[20][68] = 16'h0029;
        rom[20][69] = 16'h0011;
        rom[20][70] = 16'hFFD2;
        rom[20][71] = 16'hFFDC;
        rom[20][72] = 16'h0041;
        rom[20][73] = 16'hFFF3;
        rom[20][74] = 16'h0025;
        rom[20][75] = 16'h0018;
        rom[20][76] = 16'hFFD2;
        rom[20][77] = 16'h0000;
        rom[20][78] = 16'h000C;
        rom[20][79] = 16'h000F;
        rom[20][80] = 16'h001D;
        rom[20][81] = 16'hFFEE;
        rom[20][82] = 16'hFFEF;
        rom[20][83] = 16'h000D;
        rom[20][84] = 16'hFFD5;
        rom[20][85] = 16'h0010;
        rom[20][86] = 16'hFFF8;
        rom[20][87] = 16'h000B;
        rom[20][88] = 16'h000F;
        rom[20][89] = 16'h0015;
        rom[20][90] = 16'hFFE8;
        rom[20][91] = 16'h0004;
        rom[20][92] = 16'hFFEF;
        rom[20][93] = 16'h0019;
        rom[20][94] = 16'h0025;
        rom[20][95] = 16'hFFDB;
        rom[20][96] = 16'h000D;
        rom[20][97] = 16'h0005;
        rom[20][98] = 16'h003B;
        rom[20][99] = 16'hFFE1;
        rom[20][100] = 16'hFFF3;
        rom[20][101] = 16'hFFD4;
        rom[20][102] = 16'hFFF3;
        rom[20][103] = 16'hFFF6;
        rom[20][104] = 16'h0009;
        rom[20][105] = 16'h0014;
        rom[20][106] = 16'h0001;
        rom[20][107] = 16'hFFE7;
        rom[20][108] = 16'h0004;
        rom[20][109] = 16'h0011;
        rom[20][110] = 16'hFFD9;
        rom[20][111] = 16'h0005;
        rom[20][112] = 16'hFFE3;
        rom[20][113] = 16'hFFEB;
        rom[20][114] = 16'h000A;
        rom[20][115] = 16'hFFA1;
        rom[20][116] = 16'hFFBD;
        rom[20][117] = 16'hFFEF;
        rom[20][118] = 16'hFFF8;
        rom[20][119] = 16'hFFE4;
        rom[20][120] = 16'h0006;
        rom[20][121] = 16'h0011;
        rom[20][122] = 16'hFFA2;
        rom[20][123] = 16'hFFD7;
        rom[20][124] = 16'hFFEB;
        rom[20][125] = 16'h0019;
        rom[20][126] = 16'hFFD0;
        rom[20][127] = 16'hFFFA;
        rom[21][0] = 16'h0009;
        rom[21][1] = 16'hFFF9;
        rom[21][2] = 16'h0026;
        rom[21][3] = 16'hFFE5;
        rom[21][4] = 16'hFFCB;
        rom[21][5] = 16'h000A;
        rom[21][6] = 16'h0026;
        rom[21][7] = 16'hFFE7;
        rom[21][8] = 16'hFFDC;
        rom[21][9] = 16'h0011;
        rom[21][10] = 16'hFFCA;
        rom[21][11] = 16'hFFF2;
        rom[21][12] = 16'hFFEF;
        rom[21][13] = 16'h0006;
        rom[21][14] = 16'hFFDC;
        rom[21][15] = 16'h000E;
        rom[21][16] = 16'h0008;
        rom[21][17] = 16'hFFFD;
        rom[21][18] = 16'hFFE5;
        rom[21][19] = 16'hFFDF;
        rom[21][20] = 16'h0007;
        rom[21][21] = 16'h0007;
        rom[21][22] = 16'hFFE6;
        rom[21][23] = 16'hFFC4;
        rom[21][24] = 16'h0012;
        rom[21][25] = 16'hFFD5;
        rom[21][26] = 16'hFFD7;
        rom[21][27] = 16'hFFE6;
        rom[21][28] = 16'hFFE4;
        rom[21][29] = 16'h0025;
        rom[21][30] = 16'hFFC4;
        rom[21][31] = 16'h0028;
        rom[21][32] = 16'hFFFB;
        rom[21][33] = 16'hFFD1;
        rom[21][34] = 16'h0007;
        rom[21][35] = 16'h0032;
        rom[21][36] = 16'h0005;
        rom[21][37] = 16'hFFFE;
        rom[21][38] = 16'h0013;
        rom[21][39] = 16'h000E;
        rom[21][40] = 16'h0001;
        rom[21][41] = 16'h0009;
        rom[21][42] = 16'hFFC3;
        rom[21][43] = 16'hFFEB;
        rom[21][44] = 16'hFFF9;
        rom[21][45] = 16'h0033;
        rom[21][46] = 16'h0002;
        rom[21][47] = 16'h0009;
        rom[21][48] = 16'h001B;
        rom[21][49] = 16'h0002;
        rom[21][50] = 16'h0012;
        rom[21][51] = 16'hFFD2;
        rom[21][52] = 16'h0009;
        rom[21][53] = 16'h0001;
        rom[21][54] = 16'hFFD8;
        rom[21][55] = 16'hFFF9;
        rom[21][56] = 16'hFFFF;
        rom[21][57] = 16'hFFF4;
        rom[21][58] = 16'h0004;
        rom[21][59] = 16'hFFC8;
        rom[21][60] = 16'h0002;
        rom[21][61] = 16'h000C;
        rom[21][62] = 16'h003E;
        rom[21][63] = 16'hFFD9;
        rom[21][64] = 16'h0029;
        rom[21][65] = 16'h0016;
        rom[21][66] = 16'h0008;
        rom[21][67] = 16'hFFF8;
        rom[21][68] = 16'h001B;
        rom[21][69] = 16'hFFE6;
        rom[21][70] = 16'h0027;
        rom[21][71] = 16'h0009;
        rom[21][72] = 16'h0006;
        rom[21][73] = 16'hFFD7;
        rom[21][74] = 16'h0022;
        rom[21][75] = 16'h0000;
        rom[21][76] = 16'h0021;
        rom[21][77] = 16'hFFBE;
        rom[21][78] = 16'hFFF3;
        rom[21][79] = 16'hFFC9;
        rom[21][80] = 16'h002F;
        rom[21][81] = 16'hFFD7;
        rom[21][82] = 16'hFFF1;
        rom[21][83] = 16'hFFEC;
        rom[21][84] = 16'h0008;
        rom[21][85] = 16'h0008;
        rom[21][86] = 16'h0034;
        rom[21][87] = 16'h0001;
        rom[21][88] = 16'h000C;
        rom[21][89] = 16'h000B;
        rom[21][90] = 16'hFFF7;
        rom[21][91] = 16'h000F;
        rom[21][92] = 16'h0026;
        rom[21][93] = 16'hFFD7;
        rom[21][94] = 16'h002D;
        rom[21][95] = 16'hFFDF;
        rom[21][96] = 16'hFFD8;
        rom[21][97] = 16'h0032;
        rom[21][98] = 16'hFFF9;
        rom[21][99] = 16'hFFDA;
        rom[21][100] = 16'h0011;
        rom[21][101] = 16'h0023;
        rom[21][102] = 16'hFFEA;
        rom[21][103] = 16'hFFE4;
        rom[21][104] = 16'h0004;
        rom[21][105] = 16'hFFC8;
        rom[21][106] = 16'h002C;
        rom[21][107] = 16'hFFF0;
        rom[21][108] = 16'h001D;
        rom[21][109] = 16'hFFF9;
        rom[21][110] = 16'hFFE1;
        rom[21][111] = 16'hFFE1;
        rom[21][112] = 16'hFFD8;
        rom[21][113] = 16'hFFF7;
        rom[21][114] = 16'h0012;
        rom[21][115] = 16'h0008;
        rom[21][116] = 16'hFFBC;
        rom[21][117] = 16'h0018;
        rom[21][118] = 16'h001B;
        rom[21][119] = 16'h001B;
        rom[21][120] = 16'h001C;
        rom[21][121] = 16'hFFDC;
        rom[21][122] = 16'h001B;
        rom[21][123] = 16'hFFEF;
        rom[21][124] = 16'hFFF4;
        rom[21][125] = 16'hFFE1;
        rom[21][126] = 16'hFFF8;
        rom[21][127] = 16'hFFFD;
        rom[22][0] = 16'hFFF9;
        rom[22][1] = 16'hFFD7;
        rom[22][2] = 16'hFFD7;
        rom[22][3] = 16'h000A;
        rom[22][4] = 16'h0002;
        rom[22][5] = 16'hFFF0;
        rom[22][6] = 16'h0018;
        rom[22][7] = 16'hFFF9;
        rom[22][8] = 16'h0006;
        rom[22][9] = 16'h002C;
        rom[22][10] = 16'h0012;
        rom[22][11] = 16'hFFEE;
        rom[22][12] = 16'hFFE5;
        rom[22][13] = 16'hFFEE;
        rom[22][14] = 16'h000C;
        rom[22][15] = 16'hFFE2;
        rom[22][16] = 16'hFFD9;
        rom[22][17] = 16'hFFE3;
        rom[22][18] = 16'h0033;
        rom[22][19] = 16'hFFD1;
        rom[22][20] = 16'hFFE8;
        rom[22][21] = 16'h002D;
        rom[22][22] = 16'h001B;
        rom[22][23] = 16'h0000;
        rom[22][24] = 16'h0009;
        rom[22][25] = 16'h000D;
        rom[22][26] = 16'h0008;
        rom[22][27] = 16'h0009;
        rom[22][28] = 16'hFFD6;
        rom[22][29] = 16'hFFFC;
        rom[22][30] = 16'h002E;
        rom[22][31] = 16'h0007;
        rom[22][32] = 16'hFFD2;
        rom[22][33] = 16'h0008;
        rom[22][34] = 16'h0030;
        rom[22][35] = 16'h0013;
        rom[22][36] = 16'hFFEF;
        rom[22][37] = 16'hFFFF;
        rom[22][38] = 16'h0002;
        rom[22][39] = 16'h0002;
        rom[22][40] = 16'h000F;
        rom[22][41] = 16'h0019;
        rom[22][42] = 16'h0011;
        rom[22][43] = 16'h0003;
        rom[22][44] = 16'h002F;
        rom[22][45] = 16'h0027;
        rom[22][46] = 16'hFFE9;
        rom[22][47] = 16'hFFCE;
        rom[22][48] = 16'h0007;
        rom[22][49] = 16'h0014;
        rom[22][50] = 16'hFFDA;
        rom[22][51] = 16'h0007;
        rom[22][52] = 16'h000E;
        rom[22][53] = 16'h001F;
        rom[22][54] = 16'hFFD5;
        rom[22][55] = 16'h0037;
        rom[22][56] = 16'hFFE5;
        rom[22][57] = 16'hFFE5;
        rom[22][58] = 16'h0005;
        rom[22][59] = 16'hFFE7;
        rom[22][60] = 16'h0001;
        rom[22][61] = 16'hFFDB;
        rom[22][62] = 16'hFFFE;
        rom[22][63] = 16'hFFFC;
        rom[22][64] = 16'hFFEF;
        rom[22][65] = 16'h0002;
        rom[22][66] = 16'hFFED;
        rom[22][67] = 16'hFFDD;
        rom[22][68] = 16'h000F;
        rom[22][69] = 16'h0024;
        rom[22][70] = 16'h0022;
        rom[22][71] = 16'h0033;
        rom[22][72] = 16'h0016;
        rom[22][73] = 16'hFFE9;
        rom[22][74] = 16'hFFF1;
        rom[22][75] = 16'h001A;
        rom[22][76] = 16'hFFD0;
        rom[22][77] = 16'h0000;
        rom[22][78] = 16'hFFD4;
        rom[22][79] = 16'h0013;
        rom[22][80] = 16'h000E;
        rom[22][81] = 16'hFFAD;
        rom[22][82] = 16'hFFB3;
        rom[22][83] = 16'h000A;
        rom[22][84] = 16'hFFA6;
        rom[22][85] = 16'hFFBF;
        rom[22][86] = 16'h0011;
        rom[22][87] = 16'h0014;
        rom[22][88] = 16'h0016;
        rom[22][89] = 16'h0007;
        rom[22][90] = 16'hFFD0;
        rom[22][91] = 16'hFFE5;
        rom[22][92] = 16'h0002;
        rom[22][93] = 16'h0026;
        rom[22][94] = 16'h0026;
        rom[22][95] = 16'h001B;
        rom[22][96] = 16'h001D;
        rom[22][97] = 16'h0034;
        rom[22][98] = 16'hFFFA;
        rom[22][99] = 16'hFFE5;
        rom[22][100] = 16'h0013;
        rom[22][101] = 16'hFFF4;
        rom[22][102] = 16'hFFFE;
        rom[22][103] = 16'h0038;
        rom[22][104] = 16'h001E;
        rom[22][105] = 16'hFFDE;
        rom[22][106] = 16'hFFCD;
        rom[22][107] = 16'h0024;
        rom[22][108] = 16'hFFE4;
        rom[22][109] = 16'h0010;
        rom[22][110] = 16'hFFE1;
        rom[22][111] = 16'hFFCD;
        rom[22][112] = 16'hFFA9;
        rom[22][113] = 16'hFFD7;
        rom[22][114] = 16'hFFE1;
        rom[22][115] = 16'h002A;
        rom[22][116] = 16'h0007;
        rom[22][117] = 16'h0001;
        rom[22][118] = 16'h0067;
        rom[22][119] = 16'hFFF9;
        rom[22][120] = 16'hFFCD;
        rom[22][121] = 16'hFFE6;
        rom[22][122] = 16'h0003;
        rom[22][123] = 16'hFFE1;
        rom[22][124] = 16'hFFDA;
        rom[22][125] = 16'h000D;
        rom[22][126] = 16'h0027;
        rom[22][127] = 16'h000E;
        rom[23][0] = 16'h0001;
        rom[23][1] = 16'hFFC0;
        rom[23][2] = 16'h001C;
        rom[23][3] = 16'h002F;
        rom[23][4] = 16'hFFC2;
        rom[23][5] = 16'hFFF8;
        rom[23][6] = 16'hFFA1;
        rom[23][7] = 16'hFFE8;
        rom[23][8] = 16'hFFEC;
        rom[23][9] = 16'h000D;
        rom[23][10] = 16'hFFF5;
        rom[23][11] = 16'hFFF9;
        rom[23][12] = 16'h0001;
        rom[23][13] = 16'h0000;
        rom[23][14] = 16'h0048;
        rom[23][15] = 16'h0002;
        rom[23][16] = 16'h0016;
        rom[23][17] = 16'h0011;
        rom[23][18] = 16'h001B;
        rom[23][19] = 16'h001B;
        rom[23][20] = 16'h0002;
        rom[23][21] = 16'h0001;
        rom[23][22] = 16'hFFEF;
        rom[23][23] = 16'hFFC8;
        rom[23][24] = 16'hFFED;
        rom[23][25] = 16'h002B;
        rom[23][26] = 16'h0016;
        rom[23][27] = 16'h0026;
        rom[23][28] = 16'h001F;
        rom[23][29] = 16'h001B;
        rom[23][30] = 16'h0015;
        rom[23][31] = 16'hFFE1;
        rom[23][32] = 16'h0004;
        rom[23][33] = 16'h0016;
        rom[23][34] = 16'hFFF0;
        rom[23][35] = 16'hFFFA;
        rom[23][36] = 16'hFFD6;
        rom[23][37] = 16'hFFCA;
        rom[23][38] = 16'hFFEA;
        rom[23][39] = 16'hFFD4;
        rom[23][40] = 16'hFFE6;
        rom[23][41] = 16'hFFFC;
        rom[23][42] = 16'h001F;
        rom[23][43] = 16'h0010;
        rom[23][44] = 16'hFFFA;
        rom[23][45] = 16'h0002;
        rom[23][46] = 16'hFFFB;
        rom[23][47] = 16'hFFB8;
        rom[23][48] = 16'hFFFF;
        rom[23][49] = 16'hFFFD;
        rom[23][50] = 16'h0005;
        rom[23][51] = 16'hFFEA;
        rom[23][52] = 16'h0006;
        rom[23][53] = 16'h0014;
        rom[23][54] = 16'h0016;
        rom[23][55] = 16'hFFC1;
        rom[23][56] = 16'hFFFD;
        rom[23][57] = 16'hFFD2;
        rom[23][58] = 16'h0038;
        rom[23][59] = 16'h0015;
        rom[23][60] = 16'hFFF7;
        rom[23][61] = 16'hFFF6;
        rom[23][62] = 16'hFFE1;
        rom[23][63] = 16'hFFE8;
        rom[23][64] = 16'hFFF4;
        rom[23][65] = 16'hFFE5;
        rom[23][66] = 16'hFFA3;
        rom[23][67] = 16'hFFD8;
        rom[23][68] = 16'hFFE9;
        rom[23][69] = 16'hFFEF;
        rom[23][70] = 16'hFFED;
        rom[23][71] = 16'h0016;
        rom[23][72] = 16'h0008;
        rom[23][73] = 16'hFFDF;
        rom[23][74] = 16'h0016;
        rom[23][75] = 16'h0013;
        rom[23][76] = 16'hFFE7;
        rom[23][77] = 16'h001B;
        rom[23][78] = 16'hFFFB;
        rom[23][79] = 16'h0023;
        rom[23][80] = 16'h001E;
        rom[23][81] = 16'hFFBB;
        rom[23][82] = 16'hFFE7;
        rom[23][83] = 16'h000C;
        rom[23][84] = 16'hFFF4;
        rom[23][85] = 16'h0014;
        rom[23][86] = 16'h0016;
        rom[23][87] = 16'hFFE1;
        rom[23][88] = 16'h0004;
        rom[23][89] = 16'h000E;
        rom[23][90] = 16'h0012;
        rom[23][91] = 16'h0016;
        rom[23][92] = 16'hFFEB;
        rom[23][93] = 16'hFFE5;
        rom[23][94] = 16'h001F;
        rom[23][95] = 16'hFFE1;
        rom[23][96] = 16'hFFE1;
        rom[23][97] = 16'hFFEC;
        rom[23][98] = 16'hFFF9;
        rom[23][99] = 16'hFFAD;
        rom[23][100] = 16'hFFD4;
        rom[23][101] = 16'hFFEF;
        rom[23][102] = 16'hFFD7;
        rom[23][103] = 16'hFFD8;
        rom[23][104] = 16'hFFFE;
        rom[23][105] = 16'hFFFC;
        rom[23][106] = 16'hFFDE;
        rom[23][107] = 16'hFFFC;
        rom[23][108] = 16'h002A;
        rom[23][109] = 16'hFFF8;
        rom[23][110] = 16'hFFEA;
        rom[23][111] = 16'hFFEE;
        rom[23][112] = 16'h0033;
        rom[23][113] = 16'h0002;
        rom[23][114] = 16'hFFEA;
        rom[23][115] = 16'hFFB2;
        rom[23][116] = 16'hFFD6;
        rom[23][117] = 16'hFFEF;
        rom[23][118] = 16'hFFD5;
        rom[23][119] = 16'hFFD4;
        rom[23][120] = 16'h0005;
        rom[23][121] = 16'hFFFF;
        rom[23][122] = 16'h0009;
        rom[23][123] = 16'hFFE3;
        rom[23][124] = 16'h0014;
        rom[23][125] = 16'hFFD8;
        rom[23][126] = 16'h0020;
        rom[23][127] = 16'hFFFC;
        rom[24][0] = 16'hFFCB;
        rom[24][1] = 16'hFFF1;
        rom[24][2] = 16'hFFD5;
        rom[24][3] = 16'h001B;
        rom[24][4] = 16'h000B;
        rom[24][5] = 16'hFFF9;
        rom[24][6] = 16'hFFEE;
        rom[24][7] = 16'hFFD2;
        rom[24][8] = 16'h000C;
        rom[24][9] = 16'hFFED;
        rom[24][10] = 16'hFFEA;
        rom[24][11] = 16'hFFC4;
        rom[24][12] = 16'h0021;
        rom[24][13] = 16'hFFF1;
        rom[24][14] = 16'h001B;
        rom[24][15] = 16'h000C;
        rom[24][16] = 16'h0000;
        rom[24][17] = 16'hFFCC;
        rom[24][18] = 16'h001B;
        rom[24][19] = 16'h0011;
        rom[24][20] = 16'h0025;
        rom[24][21] = 16'hFFE2;
        rom[24][22] = 16'h0029;
        rom[24][23] = 16'hFFE0;
        rom[24][24] = 16'hFFEA;
        rom[24][25] = 16'h001D;
        rom[24][26] = 16'h0008;
        rom[24][27] = 16'h002E;
        rom[24][28] = 16'h0016;
        rom[24][29] = 16'h001A;
        rom[24][30] = 16'hFFE1;
        rom[24][31] = 16'h0010;
        rom[24][32] = 16'hFFED;
        rom[24][33] = 16'hFFEE;
        rom[24][34] = 16'h0005;
        rom[24][35] = 16'h002D;
        rom[24][36] = 16'hFFEF;
        rom[24][37] = 16'hFFE7;
        rom[24][38] = 16'hFFC1;
        rom[24][39] = 16'hFFEE;
        rom[24][40] = 16'hFFD2;
        rom[24][41] = 16'hFFFA;
        rom[24][42] = 16'h002D;
        rom[24][43] = 16'h0012;
        rom[24][44] = 16'h0023;
        rom[24][45] = 16'h0000;
        rom[24][46] = 16'hFFFA;
        rom[24][47] = 16'h0028;
        rom[24][48] = 16'hFFC8;
        rom[24][49] = 16'hFFCB;
        rom[24][50] = 16'hFFF9;
        rom[24][51] = 16'hFFFB;
        rom[24][52] = 16'hFFB0;
        rom[24][53] = 16'hFFC8;
        rom[24][54] = 16'hFFF8;
        rom[24][55] = 16'h001C;
        rom[24][56] = 16'h0018;
        rom[24][57] = 16'h002C;
        rom[24][58] = 16'h001D;
        rom[24][59] = 16'h0004;
        rom[24][60] = 16'hFFF3;
        rom[24][61] = 16'h001D;
        rom[24][62] = 16'h0012;
        rom[24][63] = 16'hFFEF;
        rom[24][64] = 16'h0016;
        rom[24][65] = 16'hFFF3;
        rom[24][66] = 16'hFFED;
        rom[24][67] = 16'hFFFE;
        rom[24][68] = 16'hFFBA;
        rom[24][69] = 16'hFFEF;
        rom[24][70] = 16'hFFE2;
        rom[24][71] = 16'hFFB9;
        rom[24][72] = 16'h000B;
        rom[24][73] = 16'hFFF8;
        rom[24][74] = 16'hFFE3;
        rom[24][75] = 16'h0002;
        rom[24][76] = 16'hFFF4;
        rom[24][77] = 16'h003C;
        rom[24][78] = 16'hFFF1;
        rom[24][79] = 16'hFFFC;
        rom[24][80] = 16'h0022;
        rom[24][81] = 16'hFFF0;
        rom[24][82] = 16'hFFDD;
        rom[24][83] = 16'h0000;
        rom[24][84] = 16'hFFFA;
        rom[24][85] = 16'hFFFE;
        rom[24][86] = 16'hFFE8;
        rom[24][87] = 16'hFFD1;
        rom[24][88] = 16'hFFD3;
        rom[24][89] = 16'hFFF9;
        rom[24][90] = 16'hFFF4;
        rom[24][91] = 16'h0004;
        rom[24][92] = 16'h000C;
        rom[24][93] = 16'h000E;
        rom[24][94] = 16'hFFD1;
        rom[24][95] = 16'hFFF6;
        rom[24][96] = 16'hFFD7;
        rom[24][97] = 16'hFFCD;
        rom[24][98] = 16'hFFFE;
        rom[24][99] = 16'h0012;
        rom[24][100] = 16'hFFDD;
        rom[24][101] = 16'hFFEF;
        rom[24][102] = 16'hFFE0;
        rom[24][103] = 16'hFFD7;
        rom[24][104] = 16'h0016;
        rom[24][105] = 16'hFFF3;
        rom[24][106] = 16'hFFF4;
        rom[24][107] = 16'hFFF6;
        rom[24][108] = 16'hFFCE;
        rom[24][109] = 16'h0025;
        rom[24][110] = 16'hFFFF;
        rom[24][111] = 16'h0002;
        rom[24][112] = 16'hFFE5;
        rom[24][113] = 16'hFFE2;
        rom[24][114] = 16'h0010;
        rom[24][115] = 16'hFFEF;
        rom[24][116] = 16'hFFF4;
        rom[24][117] = 16'hFFE1;
        rom[24][118] = 16'hFFD8;
        rom[24][119] = 16'h0007;
        rom[24][120] = 16'hFFC0;
        rom[24][121] = 16'hFFD7;
        rom[24][122] = 16'hFFE4;
        rom[24][123] = 16'h002E;
        rom[24][124] = 16'hFFFA;
        rom[24][125] = 16'hFFFE;
        rom[24][126] = 16'h002A;
        rom[24][127] = 16'h000C;
        rom[25][0] = 16'h0024;
        rom[25][1] = 16'h0006;
        rom[25][2] = 16'h0024;
        rom[25][3] = 16'hFFD7;
        rom[25][4] = 16'h0010;
        rom[25][5] = 16'hFFE9;
        rom[25][6] = 16'hFFE0;
        rom[25][7] = 16'h0007;
        rom[25][8] = 16'h0012;
        rom[25][9] = 16'hFFF6;
        rom[25][10] = 16'hFFCA;
        rom[25][11] = 16'hFFE7;
        rom[25][12] = 16'hFFF3;
        rom[25][13] = 16'h0001;
        rom[25][14] = 16'hFFF2;
        rom[25][15] = 16'h002D;
        rom[25][16] = 16'hFFF9;
        rom[25][17] = 16'h0007;
        rom[25][18] = 16'h0002;
        rom[25][19] = 16'hFFC7;
        rom[25][20] = 16'h000C;
        rom[25][21] = 16'h0010;
        rom[25][22] = 16'hFFF7;
        rom[25][23] = 16'hFFF4;
        rom[25][24] = 16'h0000;
        rom[25][25] = 16'hFFC7;
        rom[25][26] = 16'h000B;
        rom[25][27] = 16'h0002;
        rom[25][28] = 16'hFFDC;
        rom[25][29] = 16'hFFE0;
        rom[25][30] = 16'hFFFE;
        rom[25][31] = 16'h0002;
        rom[25][32] = 16'hFFFC;
        rom[25][33] = 16'h0005;
        rom[25][34] = 16'h0017;
        rom[25][35] = 16'hFFD2;
        rom[25][36] = 16'h0007;
        rom[25][37] = 16'hFFF4;
        rom[25][38] = 16'h001B;
        rom[25][39] = 16'hFFF9;
        rom[25][40] = 16'hFFBF;
        rom[25][41] = 16'hFFF4;
        rom[25][42] = 16'hFFE1;
        rom[25][43] = 16'hFFFE;
        rom[25][44] = 16'hFFF4;
        rom[25][45] = 16'hFFCD;
        rom[25][46] = 16'h0007;
        rom[25][47] = 16'hFFED;
        rom[25][48] = 16'hFFE6;
        rom[25][49] = 16'hFFAE;
        rom[25][50] = 16'h000D;
        rom[25][51] = 16'hFFCA;
        rom[25][52] = 16'h0018;
        rom[25][53] = 16'hFFB3;
        rom[25][54] = 16'h002E;
        rom[25][55] = 16'hFFFA;
        rom[25][56] = 16'hFFF3;
        rom[25][57] = 16'hFFEF;
        rom[25][58] = 16'h001E;
        rom[25][59] = 16'hFFF8;
        rom[25][60] = 16'h0021;
        rom[25][61] = 16'hFFEF;
        rom[25][62] = 16'hFFC8;
        rom[25][63] = 16'hFFF4;
        rom[25][64] = 16'h002D;
        rom[25][65] = 16'h0013;
        rom[25][66] = 16'hFFFA;
        rom[25][67] = 16'hFFF7;
        rom[25][68] = 16'hFFF0;
        rom[25][69] = 16'hFFBA;
        rom[25][70] = 16'h001D;
        rom[25][71] = 16'h002B;
        rom[25][72] = 16'h000E;
        rom[25][73] = 16'hFFFB;
        rom[25][74] = 16'hFFE2;
        rom[25][75] = 16'h000E;
        rom[25][76] = 16'h0027;
        rom[25][77] = 16'h001E;
        rom[25][78] = 16'h000D;
        rom[25][79] = 16'h0027;
        rom[25][80] = 16'hFFDF;
        rom[25][81] = 16'h0016;
        rom[25][82] = 16'hFFF0;
        rom[25][83] = 16'hFFEA;
        rom[25][84] = 16'h001D;
        rom[25][85] = 16'h0011;
        rom[25][86] = 16'hFFF2;
        rom[25][87] = 16'h001A;
        rom[25][88] = 16'h0029;
        rom[25][89] = 16'h003D;
        rom[25][90] = 16'hFFD3;
        rom[25][91] = 16'h0002;
        rom[25][92] = 16'hFFFE;
        rom[25][93] = 16'hFFCB;
        rom[25][94] = 16'hFFF1;
        rom[25][95] = 16'hFFE2;
        rom[25][96] = 16'hFFE3;
        rom[25][97] = 16'hFFD7;
        rom[25][98] = 16'hFFD0;
        rom[25][99] = 16'h000B;
        rom[25][100] = 16'h0007;
        rom[25][101] = 16'hFFEC;
        rom[25][102] = 16'hFFBA;
        rom[25][103] = 16'hFFEB;
        rom[25][104] = 16'hFFEF;
        rom[25][105] = 16'hFFE0;
        rom[25][106] = 16'h001E;
        rom[25][107] = 16'h000C;
        rom[25][108] = 16'hFFF4;
        rom[25][109] = 16'hFFCD;
        rom[25][110] = 16'h000F;
        rom[25][111] = 16'hFFD7;
        rom[25][112] = 16'hFFCC;
        rom[25][113] = 16'h000A;
        rom[25][114] = 16'hFFDE;
        rom[25][115] = 16'h0016;
        rom[25][116] = 16'h000D;
        rom[25][117] = 16'hFFEE;
        rom[25][118] = 16'h000C;
        rom[25][119] = 16'h0020;
        rom[25][120] = 16'h001E;
        rom[25][121] = 16'hFFD3;
        rom[25][122] = 16'h0027;
        rom[25][123] = 16'h000E;
        rom[25][124] = 16'h0041;
        rom[25][125] = 16'h0021;
        rom[25][126] = 16'hFFE5;
        rom[25][127] = 16'h0011;
        rom[26][0] = 16'h0007;
        rom[26][1] = 16'h000C;
        rom[26][2] = 16'hFFEF;
        rom[26][3] = 16'h0024;
        rom[26][4] = 16'h0011;
        rom[26][5] = 16'hFFFC;
        rom[26][6] = 16'h0011;
        rom[26][7] = 16'h000B;
        rom[26][8] = 16'hFFFB;
        rom[26][9] = 16'h0003;
        rom[26][10] = 16'h0020;
        rom[26][11] = 16'hFFE6;
        rom[26][12] = 16'h0005;
        rom[26][13] = 16'hFFE0;
        rom[26][14] = 16'h0016;
        rom[26][15] = 16'h0004;
        rom[26][16] = 16'hFFF9;
        rom[26][17] = 16'h0011;
        rom[26][18] = 16'hFFF0;
        rom[26][19] = 16'hFFF1;
        rom[26][20] = 16'hFFD6;
        rom[26][21] = 16'hFFE7;
        rom[26][22] = 16'h0029;
        rom[26][23] = 16'h0019;
        rom[26][24] = 16'h000A;
        rom[26][25] = 16'hFFC6;
        rom[26][26] = 16'h000D;
        rom[26][27] = 16'hFFC9;
        rom[26][28] = 16'h0016;
        rom[26][29] = 16'hFFF8;
        rom[26][30] = 16'hFFFB;
        rom[26][31] = 16'hFFB3;
        rom[26][32] = 16'hFFDC;
        rom[26][33] = 16'h0008;
        rom[26][34] = 16'hFFE9;
        rom[26][35] = 16'h000A;
        rom[26][36] = 16'hFFFD;
        rom[26][37] = 16'h000A;
        rom[26][38] = 16'h001C;
        rom[26][39] = 16'h0015;
        rom[26][40] = 16'hFFE3;
        rom[26][41] = 16'h0012;
        rom[26][42] = 16'h0010;
        rom[26][43] = 16'hFFF7;
        rom[26][44] = 16'hFFEF;
        rom[26][45] = 16'hFFC7;
        rom[26][46] = 16'h0019;
        rom[26][47] = 16'hFFED;
        rom[26][48] = 16'hFFDC;
        rom[26][49] = 16'hFFA6;
        rom[26][50] = 16'hFFDC;
        rom[26][51] = 16'hFFF3;
        rom[26][52] = 16'h0037;
        rom[26][53] = 16'hFFC0;
        rom[26][54] = 16'hFFA2;
        rom[26][55] = 16'hFFBA;
        rom[26][56] = 16'hFFE8;
        rom[26][57] = 16'hFFEF;
        rom[26][58] = 16'h0038;
        rom[26][59] = 16'h000F;
        rom[26][60] = 16'hFFD7;
        rom[26][61] = 16'hFFCD;
        rom[26][62] = 16'h0002;
        rom[26][63] = 16'hFFF6;
        rom[26][64] = 16'h000A;
        rom[26][65] = 16'h001F;
        rom[26][66] = 16'h0007;
        rom[26][67] = 16'hFFEC;
        rom[26][68] = 16'h0012;
        rom[26][69] = 16'hFFF4;
        rom[26][70] = 16'h000B;
        rom[26][71] = 16'h0033;
        rom[26][72] = 16'hFFE8;
        rom[26][73] = 16'hFFF4;
        rom[26][74] = 16'hFFEB;
        rom[26][75] = 16'hFFF4;
        rom[26][76] = 16'h0002;
        rom[26][77] = 16'h0036;
        rom[26][78] = 16'h0025;
        rom[26][79] = 16'h0010;
        rom[26][80] = 16'hFFF9;
        rom[26][81] = 16'hFFF2;
        rom[26][82] = 16'h0024;
        rom[26][83] = 16'hFFDB;
        rom[26][84] = 16'h0027;
        rom[26][85] = 16'hFFD2;
        rom[26][86] = 16'h0005;
        rom[26][87] = 16'hFFFB;
        rom[26][88] = 16'hFFF7;
        rom[26][89] = 16'hFFDE;
        rom[26][90] = 16'h0002;
        rom[26][91] = 16'hFFEA;
        rom[26][92] = 16'hFFEB;
        rom[26][93] = 16'h0031;
        rom[26][94] = 16'hFFFE;
        rom[26][95] = 16'h0031;
        rom[26][96] = 16'h001B;
        rom[26][97] = 16'h0017;
        rom[26][98] = 16'hFFC3;
        rom[26][99] = 16'hFFEA;
        rom[26][100] = 16'h0031;
        rom[26][101] = 16'hFFF9;
        rom[26][102] = 16'hFFF0;
        rom[26][103] = 16'h0008;
        rom[26][104] = 16'hFFE9;
        rom[26][105] = 16'hFFF9;
        rom[26][106] = 16'h0033;
        rom[26][107] = 16'hFFDD;
        rom[26][108] = 16'hFFD5;
        rom[26][109] = 16'h0007;
        rom[26][110] = 16'hFFF0;
        rom[26][111] = 16'h0043;
        rom[26][112] = 16'h0002;
        rom[26][113] = 16'hFFD3;
        rom[26][114] = 16'hFFC3;
        rom[26][115] = 16'hFFCC;
        rom[26][116] = 16'h000D;
        rom[26][117] = 16'h0029;
        rom[26][118] = 16'h0007;
        rom[26][119] = 16'h0011;
        rom[26][120] = 16'hFFDA;
        rom[26][121] = 16'h0005;
        rom[26][122] = 16'hFFDA;
        rom[26][123] = 16'h0018;
        rom[26][124] = 16'hFFF4;
        rom[26][125] = 16'hFFED;
        rom[26][126] = 16'hFFFE;
        rom[26][127] = 16'h0016;
        rom[27][0] = 16'h000E;
        rom[27][1] = 16'h0017;
        rom[27][2] = 16'hFFD6;
        rom[27][3] = 16'h0013;
        rom[27][4] = 16'h0034;
        rom[27][5] = 16'h0000;
        rom[27][6] = 16'h001D;
        rom[27][7] = 16'h0007;
        rom[27][8] = 16'hFFE4;
        rom[27][9] = 16'hFFD1;
        rom[27][10] = 16'h0014;
        rom[27][11] = 16'hFFF7;
        rom[27][12] = 16'hFFF1;
        rom[27][13] = 16'h0011;
        rom[27][14] = 16'hFFE9;
        rom[27][15] = 16'hFFC5;
        rom[27][16] = 16'hFFF4;
        rom[27][17] = 16'h0002;
        rom[27][18] = 16'hFFEB;
        rom[27][19] = 16'h000A;
        rom[27][20] = 16'h001B;
        rom[27][21] = 16'h000D;
        rom[27][22] = 16'h0024;
        rom[27][23] = 16'h0010;
        rom[27][24] = 16'hFFC6;
        rom[27][25] = 16'hFFE5;
        rom[27][26] = 16'h0028;
        rom[27][27] = 16'hFFD9;
        rom[27][28] = 16'h0001;
        rom[27][29] = 16'hFFDB;
        rom[27][30] = 16'h0004;
        rom[27][31] = 16'hFFF4;
        rom[27][32] = 16'hFFFE;
        rom[27][33] = 16'hFFBD;
        rom[27][34] = 16'hFFEA;
        rom[27][35] = 16'hFFD8;
        rom[27][36] = 16'h0002;
        rom[27][37] = 16'h0026;
        rom[27][38] = 16'hFFC0;
        rom[27][39] = 16'hFFFD;
        rom[27][40] = 16'h0008;
        rom[27][41] = 16'hFFED;
        rom[27][42] = 16'h001A;
        rom[27][43] = 16'hFFD4;
        rom[27][44] = 16'hFFDC;
        rom[27][45] = 16'hFFF4;
        rom[27][46] = 16'hFFDC;
        rom[27][47] = 16'hFFDE;
        rom[27][48] = 16'hFFDC;
        rom[27][49] = 16'hFFFA;
        rom[27][50] = 16'hFFD4;
        rom[27][51] = 16'h0020;
        rom[27][52] = 16'h002D;
        rom[27][53] = 16'hFFFB;
        rom[27][54] = 16'h000A;
        rom[27][55] = 16'hFFFA;
        rom[27][56] = 16'hFFD7;
        rom[27][57] = 16'h0007;
        rom[27][58] = 16'hFFD9;
        rom[27][59] = 16'h000E;
        rom[27][60] = 16'h0002;
        rom[27][61] = 16'hFFBC;
        rom[27][62] = 16'hFFEA;
        rom[27][63] = 16'hFFF8;
        rom[27][64] = 16'h0006;
        rom[27][65] = 16'hFFEA;
        rom[27][66] = 16'h0011;
        rom[27][67] = 16'h002E;
        rom[27][68] = 16'hFFF1;
        rom[27][69] = 16'h0038;
        rom[27][70] = 16'h0002;
        rom[27][71] = 16'hFFF2;
        rom[27][72] = 16'h0004;
        rom[27][73] = 16'hFFF4;
        rom[27][74] = 16'hFFCA;
        rom[27][75] = 16'hFFC3;
        rom[27][76] = 16'h0005;
        rom[27][77] = 16'hFFF0;
        rom[27][78] = 16'h0011;
        rom[27][79] = 16'hFFE5;
        rom[27][80] = 16'hFFD1;
        rom[27][81] = 16'h0007;
        rom[27][82] = 16'h000A;
        rom[27][83] = 16'hFFEA;
        rom[27][84] = 16'hFFD9;
        rom[27][85] = 16'hFFC8;
        rom[27][86] = 16'hFFD1;
        rom[27][87] = 16'h001E;
        rom[27][88] = 16'h000B;
        rom[27][89] = 16'hFFCF;
        rom[27][90] = 16'h0010;
        rom[27][91] = 16'h002D;
        rom[27][92] = 16'hFFD7;
        rom[27][93] = 16'h0006;
        rom[27][94] = 16'hFFF5;
        rom[27][95] = 16'h0002;
        rom[27][96] = 16'hFFEE;
        rom[27][97] = 16'h0017;
        rom[27][98] = 16'h0002;
        rom[27][99] = 16'h0009;
        rom[27][100] = 16'h0016;
        rom[27][101] = 16'h003F;
        rom[27][102] = 16'h002E;
        rom[27][103] = 16'h0024;
        rom[27][104] = 16'h002D;
        rom[27][105] = 16'hFFFE;
        rom[27][106] = 16'h001F;
        rom[27][107] = 16'h0010;
        rom[27][108] = 16'h000C;
        rom[27][109] = 16'h0007;
        rom[27][110] = 16'h0002;
        rom[27][111] = 16'h001A;
        rom[27][112] = 16'h0014;
        rom[27][113] = 16'h0018;
        rom[27][114] = 16'h0019;
        rom[27][115] = 16'hFFFC;
        rom[27][116] = 16'hFFFD;
        rom[27][117] = 16'h0009;
        rom[27][118] = 16'hFFE0;
        rom[27][119] = 16'hFFE3;
        rom[27][120] = 16'h0004;
        rom[27][121] = 16'hFFEB;
        rom[27][122] = 16'hFFE9;
        rom[27][123] = 16'hFFBC;
        rom[27][124] = 16'hFFF4;
        rom[27][125] = 16'hFFF9;
        rom[27][126] = 16'h001A;
        rom[27][127] = 16'h0022;
        rom[28][0] = 16'hFFE1;
        rom[28][1] = 16'hFFF1;
        rom[28][2] = 16'hFFDE;
        rom[28][3] = 16'hFFE1;
        rom[28][4] = 16'hFFFE;
        rom[28][5] = 16'hFFD0;
        rom[28][6] = 16'hFFE9;
        rom[28][7] = 16'hFFFD;
        rom[28][8] = 16'h0003;
        rom[28][9] = 16'h0025;
        rom[28][10] = 16'h001E;
        rom[28][11] = 16'h0028;
        rom[28][12] = 16'h0023;
        rom[28][13] = 16'hFFF1;
        rom[28][14] = 16'hFFE7;
        rom[28][15] = 16'h000C;
        rom[28][16] = 16'h0002;
        rom[28][17] = 16'hFFFE;
        rom[28][18] = 16'hFFFF;
        rom[28][19] = 16'hFFBF;
        rom[28][20] = 16'h0007;
        rom[28][21] = 16'h0024;
        rom[28][22] = 16'hFFE8;
        rom[28][23] = 16'hFFDC;
        rom[28][24] = 16'h0024;
        rom[28][25] = 16'h0011;
        rom[28][26] = 16'hFFFE;
        rom[28][27] = 16'h0016;
        rom[28][28] = 16'hFFD6;
        rom[28][29] = 16'h0012;
        rom[28][30] = 16'h001E;
        rom[28][31] = 16'h0010;
        rom[28][32] = 16'h0011;
        rom[28][33] = 16'h0022;
        rom[28][34] = 16'h0001;
        rom[28][35] = 16'h002E;
        rom[28][36] = 16'h0005;
        rom[28][37] = 16'hFFDF;
        rom[28][38] = 16'h000C;
        rom[28][39] = 16'h0008;
        rom[28][40] = 16'h002A;
        rom[28][41] = 16'hFFE6;
        rom[28][42] = 16'h001A;
        rom[28][43] = 16'hFFCF;
        rom[28][44] = 16'h001B;
        rom[28][45] = 16'h002C;
        rom[28][46] = 16'h0017;
        rom[28][47] = 16'hFFEC;
        rom[28][48] = 16'h000A;
        rom[28][49] = 16'hFFED;
        rom[28][50] = 16'h0004;
        rom[28][51] = 16'hFFEF;
        rom[28][52] = 16'hFFC7;
        rom[28][53] = 16'h0011;
        rom[28][54] = 16'hFFFE;
        rom[28][55] = 16'h001D;
        rom[28][56] = 16'h0033;
        rom[28][57] = 16'hFFC8;
        rom[28][58] = 16'hFFFB;
        rom[28][59] = 16'h0022;
        rom[28][60] = 16'h001C;
        rom[28][61] = 16'hFFEF;
        rom[28][62] = 16'hFFEA;
        rom[28][63] = 16'hFFBA;
        rom[28][64] = 16'hFFE0;
        rom[28][65] = 16'h0024;
        rom[28][66] = 16'hFFEA;
        rom[28][67] = 16'hFFE7;
        rom[28][68] = 16'hFFDA;
        rom[28][69] = 16'hFFEF;
        rom[28][70] = 16'h0011;
        rom[28][71] = 16'hFFCD;
        rom[28][72] = 16'hFFEA;
        rom[28][73] = 16'h002A;
        rom[28][74] = 16'hFFE6;
        rom[28][75] = 16'h000D;
        rom[28][76] = 16'hFFFB;
        rom[28][77] = 16'h002A;
        rom[28][78] = 16'hFFBF;
        rom[28][79] = 16'h000F;
        rom[28][80] = 16'hFFBF;
        rom[28][81] = 16'hFFEA;
        rom[28][82] = 16'hFFBD;
        rom[28][83] = 16'h0032;
        rom[28][84] = 16'hFFF2;
        rom[28][85] = 16'hFFF2;
        rom[28][86] = 16'hFFF8;
        rom[28][87] = 16'hFFF7;
        rom[28][88] = 16'h0049;
        rom[28][89] = 16'h0004;
        rom[28][90] = 16'hFFDA;
        rom[28][91] = 16'hFFAA;
        rom[28][92] = 16'h001F;
        rom[28][93] = 16'h0004;
        rom[28][94] = 16'h0011;
        rom[28][95] = 16'hFFEB;
        rom[28][96] = 16'hFFEF;
        rom[28][97] = 16'hFFE1;
        rom[28][98] = 16'hFFB7;
        rom[28][99] = 16'hFFF3;
        rom[28][100] = 16'hFFE1;
        rom[28][101] = 16'hFFE8;
        rom[28][102] = 16'h0020;
        rom[28][103] = 16'hFFE6;
        rom[28][104] = 16'hFFD7;
        rom[28][105] = 16'hFFD7;
        rom[28][106] = 16'hFFDA;
        rom[28][107] = 16'hFFEF;
        rom[28][108] = 16'h0013;
        rom[28][109] = 16'h000E;
        rom[28][110] = 16'hFFEA;
        rom[28][111] = 16'hFFCE;
        rom[28][112] = 16'hFFEF;
        rom[28][113] = 16'h000A;
        rom[28][114] = 16'h0019;
        rom[28][115] = 16'h0027;
        rom[28][116] = 16'h0028;
        rom[28][117] = 16'hFFEC;
        rom[28][118] = 16'hFFB3;
        rom[28][119] = 16'h002E;
        rom[28][120] = 16'h0020;
        rom[28][121] = 16'hFFCC;
        rom[28][122] = 16'h0016;
        rom[28][123] = 16'hFFFE;
        rom[28][124] = 16'h0009;
        rom[28][125] = 16'hFFE9;
        rom[28][126] = 16'hFFB4;
        rom[28][127] = 16'hFFC6;
        rom[29][0] = 16'hFFD5;
        rom[29][1] = 16'h0000;
        rom[29][2] = 16'h0016;
        rom[29][3] = 16'hFFD4;
        rom[29][4] = 16'h000F;
        rom[29][5] = 16'h001A;
        rom[29][6] = 16'h0048;
        rom[29][7] = 16'hFFF5;
        rom[29][8] = 16'h0001;
        rom[29][9] = 16'hFFFE;
        rom[29][10] = 16'h001D;
        rom[29][11] = 16'h0005;
        rom[29][12] = 16'hFFCD;
        rom[29][13] = 16'h0001;
        rom[29][14] = 16'hFFEC;
        rom[29][15] = 16'hFFBF;
        rom[29][16] = 16'h0002;
        rom[29][17] = 16'h000B;
        rom[29][18] = 16'h0002;
        rom[29][19] = 16'hFFF8;
        rom[29][20] = 16'h0035;
        rom[29][21] = 16'hFFF0;
        rom[29][22] = 16'hFFF9;
        rom[29][23] = 16'h000F;
        rom[29][24] = 16'hFFDE;
        rom[29][25] = 16'h001C;
        rom[29][26] = 16'h002A;
        rom[29][27] = 16'h0000;
        rom[29][28] = 16'hFFC9;
        rom[29][29] = 16'hFFB4;
        rom[29][30] = 16'h0050;
        rom[29][31] = 16'hFFD7;
        rom[29][32] = 16'h001E;
        rom[29][33] = 16'hFFC7;
        rom[29][34] = 16'h0028;
        rom[29][35] = 16'hFFBE;
        rom[29][36] = 16'h0007;
        rom[29][37] = 16'h0017;
        rom[29][38] = 16'hFFDD;
        rom[29][39] = 16'hFFCD;
        rom[29][40] = 16'hFFEE;
        rom[29][41] = 16'hFFEE;
        rom[29][42] = 16'hFFEA;
        rom[29][43] = 16'hFFE9;
        rom[29][44] = 16'hFFCD;
        rom[29][45] = 16'hFFC5;
        rom[29][46] = 16'h0006;
        rom[29][47] = 16'hFFCD;
        rom[29][48] = 16'hFFE5;
        rom[29][49] = 16'h001B;
        rom[29][50] = 16'hFFDF;
        rom[29][51] = 16'h0014;
        rom[29][52] = 16'hFFFF;
        rom[29][53] = 16'hFFC5;
        rom[29][54] = 16'hFFFE;
        rom[29][55] = 16'hFFFC;
        rom[29][56] = 16'hFFFE;
        rom[29][57] = 16'hFFE4;
        rom[29][58] = 16'hFFA3;
        rom[29][59] = 16'h001B;
        rom[29][60] = 16'hFFF4;
        rom[29][61] = 16'hFFC8;
        rom[29][62] = 16'h000D;
        rom[29][63] = 16'h0038;
        rom[29][64] = 16'hFFDB;
        rom[29][65] = 16'hFFD0;
        rom[29][66] = 16'h001D;
        rom[29][67] = 16'h0019;
        rom[29][68] = 16'hFFD4;
        rom[29][69] = 16'hFFCD;
        rom[29][70] = 16'hFFCC;
        rom[29][71] = 16'h0019;
        rom[29][72] = 16'h0011;
        rom[29][73] = 16'h0006;
        rom[29][74] = 16'hFFD2;
        rom[29][75] = 16'hFFF5;
        rom[29][76] = 16'h001F;
        rom[29][77] = 16'h000C;
        rom[29][78] = 16'hFFEC;
        rom[29][79] = 16'hFFE7;
        rom[29][80] = 16'hFFD9;
        rom[29][81] = 16'hFFD7;
        rom[29][82] = 16'h0023;
        rom[29][83] = 16'hFFD3;
        rom[29][84] = 16'hFFCD;
        rom[29][85] = 16'hFFEA;
        rom[29][86] = 16'h0015;
        rom[29][87] = 16'h000D;
        rom[29][88] = 16'h0007;
        rom[29][89] = 16'hFFBF;
        rom[29][90] = 16'h0011;
        rom[29][91] = 16'h000A;
        rom[29][92] = 16'h0009;
        rom[29][93] = 16'hFFC8;
        rom[29][94] = 16'hFFCB;
        rom[29][95] = 16'hFFB2;
        rom[29][96] = 16'hFFDF;
        rom[29][97] = 16'h002F;
        rom[29][98] = 16'h0038;
        rom[29][99] = 16'h000C;
        rom[29][100] = 16'h001E;
        rom[29][101] = 16'hFFEF;
        rom[29][102] = 16'h0029;
        rom[29][103] = 16'h0005;
        rom[29][104] = 16'hFFE1;
        rom[29][105] = 16'hFFDD;
        rom[29][106] = 16'h001E;
        rom[29][107] = 16'hFFE2;
        rom[29][108] = 16'h0019;
        rom[29][109] = 16'hFFA3;
        rom[29][110] = 16'hFFF8;
        rom[29][111] = 16'hFFF0;
        rom[29][112] = 16'hFFEF;
        rom[29][113] = 16'hFFFB;
        rom[29][114] = 16'h000D;
        rom[29][115] = 16'h002D;
        rom[29][116] = 16'h0018;
        rom[29][117] = 16'h0003;
        rom[29][118] = 16'h0015;
        rom[29][119] = 16'hFFBC;
        rom[29][120] = 16'h0012;
        rom[29][121] = 16'h0011;
        rom[29][122] = 16'h0016;
        rom[29][123] = 16'h0000;
        rom[29][124] = 16'hFFF6;
        rom[29][125] = 16'hFFD2;
        rom[29][126] = 16'h0002;
        rom[29][127] = 16'h0023;
        rom[30][0] = 16'hFFFE;
        rom[30][1] = 16'hFFE1;
        rom[30][2] = 16'hFFE8;
        rom[30][3] = 16'h0007;
        rom[30][4] = 16'hFFE1;
        rom[30][5] = 16'h0014;
        rom[30][6] = 16'hFFE0;
        rom[30][7] = 16'hFFFC;
        rom[30][8] = 16'hFFEF;
        rom[30][9] = 16'hFFF7;
        rom[30][10] = 16'h0028;
        rom[30][11] = 16'hFFB3;
        rom[30][12] = 16'h0022;
        rom[30][13] = 16'h0017;
        rom[30][14] = 16'hFFEF;
        rom[30][15] = 16'h0029;
        rom[30][16] = 16'hFFF2;
        rom[30][17] = 16'h0007;
        rom[30][18] = 16'hFFEC;
        rom[30][19] = 16'h0016;
        rom[30][20] = 16'hFFD4;
        rom[30][21] = 16'h0007;
        rom[30][22] = 16'hFFE9;
        rom[30][23] = 16'hFFF7;
        rom[30][24] = 16'h0027;
        rom[30][25] = 16'hFFB0;
        rom[30][26] = 16'h0010;
        rom[30][27] = 16'hFFC1;
        rom[30][28] = 16'h0026;
        rom[30][29] = 16'h0014;
        rom[30][30] = 16'h0020;
        rom[30][31] = 16'hFFEE;
        rom[30][32] = 16'hFFDB;
        rom[30][33] = 16'h0028;
        rom[30][34] = 16'hFFC4;
        rom[30][35] = 16'hFFFC;
        rom[30][36] = 16'hFFEF;
        rom[30][37] = 16'hFFF8;
        rom[30][38] = 16'hFFC4;
        rom[30][39] = 16'h0026;
        rom[30][40] = 16'h001F;
        rom[30][41] = 16'h0006;
        rom[30][42] = 16'h0007;
        rom[30][43] = 16'hFFE6;
        rom[30][44] = 16'h001A;
        rom[30][45] = 16'hFFCA;
        rom[30][46] = 16'hFFDD;
        rom[30][47] = 16'h0003;
        rom[30][48] = 16'hFFEF;
        rom[30][49] = 16'h000D;
        rom[30][50] = 16'hFFDB;
        rom[30][51] = 16'h000F;
        rom[30][52] = 16'hFFB2;
        rom[30][53] = 16'h0020;
        rom[30][54] = 16'h0002;
        rom[30][55] = 16'hFFF9;
        rom[30][56] = 16'h002D;
        rom[30][57] = 16'h0011;
        rom[30][58] = 16'hFFF9;
        rom[30][59] = 16'hFFF0;
        rom[30][60] = 16'h003F;
        rom[30][61] = 16'h000C;
        rom[30][62] = 16'hFFC2;
        rom[30][63] = 16'hFFE1;
        rom[30][64] = 16'h001D;
        rom[30][65] = 16'hFFCD;
        rom[30][66] = 16'hFFFE;
        rom[30][67] = 16'h000F;
        rom[30][68] = 16'h000A;
        rom[30][69] = 16'h0012;
        rom[30][70] = 16'hFFE8;
        rom[30][71] = 16'hFFDD;
        rom[30][72] = 16'hFFF7;
        rom[30][73] = 16'h000A;
        rom[30][74] = 16'hFFFB;
        rom[30][75] = 16'h000A;
        rom[30][76] = 16'hFFFB;
        rom[30][77] = 16'h0019;
        rom[30][78] = 16'h001A;
        rom[30][79] = 16'h0003;
        rom[30][80] = 16'hFFFA;
        rom[30][81] = 16'hFFF6;
        rom[30][82] = 16'h0005;
        rom[30][83] = 16'h0013;
        rom[30][84] = 16'hFFD7;
        rom[30][85] = 16'h0019;
        rom[30][86] = 16'h001E;
        rom[30][87] = 16'hFFC6;
        rom[30][88] = 16'hFFB0;
        rom[30][89] = 16'h0007;
        rom[30][90] = 16'hFFF8;
        rom[30][91] = 16'h0004;
        rom[30][92] = 16'hFFBB;
        rom[30][93] = 16'hFFED;
        rom[30][94] = 16'h0016;
        rom[30][95] = 16'hFFE1;
        rom[30][96] = 16'h0007;
        rom[30][97] = 16'h0024;
        rom[30][98] = 16'h0011;
        rom[30][99] = 16'h0009;
        rom[30][100] = 16'h0033;
        rom[30][101] = 16'hFFFA;
        rom[30][102] = 16'hFFF4;
        rom[30][103] = 16'hFFC3;
        rom[30][104] = 16'h0000;
        rom[30][105] = 16'hFF99;
        rom[30][106] = 16'h0024;
        rom[30][107] = 16'hFFD4;
        rom[30][108] = 16'h0010;
        rom[30][109] = 16'hFFF0;
        rom[30][110] = 16'h000D;
        rom[30][111] = 16'hFFFA;
        rom[30][112] = 16'h0021;
        rom[30][113] = 16'h000A;
        rom[30][114] = 16'hFFEB;
        rom[30][115] = 16'hFFCF;
        rom[30][116] = 16'hFFB2;
        rom[30][117] = 16'h0010;
        rom[30][118] = 16'h001E;
        rom[30][119] = 16'hFFDB;
        rom[30][120] = 16'h002C;
        rom[30][121] = 16'h001E;
        rom[30][122] = 16'hFFBF;
        rom[30][123] = 16'hFFCF;
        rom[30][124] = 16'hFFF2;
        rom[30][125] = 16'hFFFD;
        rom[30][126] = 16'hFFDB;
        rom[30][127] = 16'hFFE1;
        rom[31][0] = 16'hFFFB;
        rom[31][1] = 16'h000C;
        rom[31][2] = 16'h0025;
        rom[31][3] = 16'hFFDC;
        rom[31][4] = 16'hFFEE;
        rom[31][5] = 16'h002E;
        rom[31][6] = 16'h0007;
        rom[31][7] = 16'h000C;
        rom[31][8] = 16'h0002;
        rom[31][9] = 16'h0029;
        rom[31][10] = 16'h0033;
        rom[31][11] = 16'hFFE2;
        rom[31][12] = 16'h0001;
        rom[31][13] = 16'hFFC1;
        rom[31][14] = 16'h0066;
        rom[31][15] = 16'h0011;
        rom[31][16] = 16'hFFA4;
        rom[31][17] = 16'hFFC4;
        rom[31][18] = 16'h002B;
        rom[31][19] = 16'hFFD7;
        rom[31][20] = 16'h0017;
        rom[31][21] = 16'h0014;
        rom[31][22] = 16'h001F;
        rom[31][23] = 16'h0007;
        rom[31][24] = 16'h0015;
        rom[31][25] = 16'h0018;
        rom[31][26] = 16'hFFF4;
        rom[31][27] = 16'hFFD6;
        rom[31][28] = 16'hFFD1;
        rom[31][29] = 16'hFFD0;
        rom[31][30] = 16'h0007;
        rom[31][31] = 16'hFFD6;
        rom[31][32] = 16'h000A;
        rom[31][33] = 16'hFFF6;
        rom[31][34] = 16'hFFDF;
        rom[31][35] = 16'hFFDE;
        rom[31][36] = 16'hFFFE;
        rom[31][37] = 16'h0022;
        rom[31][38] = 16'h0029;
        rom[31][39] = 16'hFFE5;
        rom[31][40] = 16'hFFCA;
        rom[31][41] = 16'h0034;
        rom[31][42] = 16'h000C;
        rom[31][43] = 16'h0011;
        rom[31][44] = 16'hFFCC;
        rom[31][45] = 16'h0004;
        rom[31][46] = 16'h001B;
        rom[31][47] = 16'h0024;
        rom[31][48] = 16'hFFE2;
        rom[31][49] = 16'h000E;
        rom[31][50] = 16'h0002;
        rom[31][51] = 16'hFFC0;
        rom[31][52] = 16'h0018;
        rom[31][53] = 16'hFFCA;
        rom[31][54] = 16'h0000;
        rom[31][55] = 16'h003F;
        rom[31][56] = 16'hFFFB;
        rom[31][57] = 16'hFFC3;
        rom[31][58] = 16'hFFE8;
        rom[31][59] = 16'h002C;
        rom[31][60] = 16'hFFE5;
        rom[31][61] = 16'h000A;
        rom[31][62] = 16'h002F;
        rom[31][63] = 16'h0011;
        rom[31][64] = 16'hFFFB;
        rom[31][65] = 16'hFFDC;
        rom[31][66] = 16'h0027;
        rom[31][67] = 16'h0010;
        rom[31][68] = 16'hFFE3;
        rom[31][69] = 16'h001B;
        rom[31][70] = 16'h0012;
        rom[31][71] = 16'hFFDC;
        rom[31][72] = 16'hFFB7;
        rom[31][73] = 16'hFFF2;
        rom[31][74] = 16'hFFE1;
        rom[31][75] = 16'h002F;
        rom[31][76] = 16'hFFDE;
        rom[31][77] = 16'hFFD7;
        rom[31][78] = 16'h001B;
        rom[31][79] = 16'hFFF7;
        rom[31][80] = 16'h001E;
        rom[31][81] = 16'hFFFB;
        rom[31][82] = 16'h0011;
        rom[31][83] = 16'h0008;
        rom[31][84] = 16'hFFEA;
        rom[31][85] = 16'h0003;
        rom[31][86] = 16'hFFD3;
        rom[31][87] = 16'hFFE7;
        rom[31][88] = 16'hFFFB;
        rom[31][89] = 16'hFFE5;
        rom[31][90] = 16'h002E;
        rom[31][91] = 16'hFFC1;
        rom[31][92] = 16'hFFF4;
        rom[31][93] = 16'hFFEA;
        rom[31][94] = 16'hFFD6;
        rom[31][95] = 16'hFFF4;
        rom[31][96] = 16'hFFF3;
        rom[31][97] = 16'hFFD6;
        rom[31][98] = 16'hFFA9;
        rom[31][99] = 16'hFFF3;
        rom[31][100] = 16'hFFFA;
        rom[31][101] = 16'h0019;
        rom[31][102] = 16'hFFFE;
        rom[31][103] = 16'hFFF6;
        rom[31][104] = 16'hFFE8;
        rom[31][105] = 16'hFFFC;
        rom[31][106] = 16'hFFD5;
        rom[31][107] = 16'h002A;
        rom[31][108] = 16'hFFEF;
        rom[31][109] = 16'hFFE1;
        rom[31][110] = 16'hFFFA;
        rom[31][111] = 16'h0001;
        rom[31][112] = 16'hFFEF;
        rom[31][113] = 16'h002D;
        rom[31][114] = 16'hFFD2;
        rom[31][115] = 16'hFFFB;
        rom[31][116] = 16'hFFF9;
        rom[31][117] = 16'h0026;
        rom[31][118] = 16'h0024;
        rom[31][119] = 16'h0031;
        rom[31][120] = 16'hFFF7;
        rom[31][121] = 16'h0011;
        rom[31][122] = 16'hFFF4;
        rom[31][123] = 16'hFFE3;
        rom[31][124] = 16'hFFE5;
        rom[31][125] = 16'h000B;
        rom[31][126] = 16'hFFC2;
        rom[31][127] = 16'h001B;
        rom[32][0] = 16'hFFEB;
        rom[32][1] = 16'h0022;
        rom[32][2] = 16'hFFEE;
        rom[32][3] = 16'hFFF7;
        rom[32][4] = 16'h0011;
        rom[32][5] = 16'h000D;
        rom[32][6] = 16'h0013;
        rom[32][7] = 16'h0010;
        rom[32][8] = 16'hFFEF;
        rom[32][9] = 16'h0002;
        rom[32][10] = 16'hFFDA;
        rom[32][11] = 16'h001D;
        rom[32][12] = 16'h0000;
        rom[32][13] = 16'hFFF1;
        rom[32][14] = 16'h0000;
        rom[32][15] = 16'hFFED;
        rom[32][16] = 16'h0039;
        rom[32][17] = 16'h0018;
        rom[32][18] = 16'hFFF3;
        rom[32][19] = 16'hFFFD;
        rom[32][20] = 16'h0000;
        rom[32][21] = 16'hFFF3;
        rom[32][22] = 16'hFFFB;
        rom[32][23] = 16'hFFFE;
        rom[32][24] = 16'hFFF8;
        rom[32][25] = 16'hFFEF;
        rom[32][26] = 16'h0023;
        rom[32][27] = 16'hFFF4;
        rom[32][28] = 16'hFFFE;
        rom[32][29] = 16'hFFD3;
        rom[32][30] = 16'h0016;
        rom[32][31] = 16'hFFE7;
        rom[32][32] = 16'hFFC8;
        rom[32][33] = 16'hFFFF;
        rom[32][34] = 16'hFFF1;
        rom[32][35] = 16'hFFD8;
        rom[32][36] = 16'h0007;
        rom[32][37] = 16'h0007;
        rom[32][38] = 16'hFFF6;
        rom[32][39] = 16'hFFAB;
        rom[32][40] = 16'hFFEF;
        rom[32][41] = 16'hFFE0;
        rom[32][42] = 16'h0014;
        rom[32][43] = 16'hFFEF;
        rom[32][44] = 16'hFFE9;
        rom[32][45] = 16'hFFB1;
        rom[32][46] = 16'h0020;
        rom[32][47] = 16'h0007;
        rom[32][48] = 16'h0016;
        rom[32][49] = 16'hFFEB;
        rom[32][50] = 16'h0014;
        rom[32][51] = 16'h000C;
        rom[32][52] = 16'hFFEC;
        rom[32][53] = 16'hFFE9;
        rom[32][54] = 16'hFFF9;
        rom[32][55] = 16'hFFDB;
        rom[32][56] = 16'h000A;
        rom[32][57] = 16'h0007;
        rom[32][58] = 16'h0013;
        rom[32][59] = 16'h000D;
        rom[32][60] = 16'hFFFF;
        rom[32][61] = 16'hFFF3;
        rom[32][62] = 16'hFFD0;
        rom[32][63] = 16'h0018;
        rom[32][64] = 16'hFFFD;
        rom[32][65] = 16'hFFE7;
        rom[32][66] = 16'h001B;
        rom[32][67] = 16'h0007;
        rom[32][68] = 16'hFFFC;
        rom[32][69] = 16'hFFE1;
        rom[32][70] = 16'hFFD7;
        rom[32][71] = 16'hFFE9;
        rom[32][72] = 16'hFFEA;
        rom[32][73] = 16'h000C;
        rom[32][74] = 16'h0007;
        rom[32][75] = 16'h0016;
        rom[32][76] = 16'h002A;
        rom[32][77] = 16'h000B;
        rom[32][78] = 16'hFFCA;
        rom[32][79] = 16'hFFF5;
        rom[32][80] = 16'h000D;
        rom[32][81] = 16'h0013;
        rom[32][82] = 16'h0011;
        rom[32][83] = 16'hFFC8;
        rom[32][84] = 16'h0010;
        rom[32][85] = 16'h0029;
        rom[32][86] = 16'hFFE5;
        rom[32][87] = 16'h002A;
        rom[32][88] = 16'hFFBF;
        rom[32][89] = 16'hFFD5;
        rom[32][90] = 16'h0002;
        rom[32][91] = 16'h001B;
        rom[32][92] = 16'h0021;
        rom[32][93] = 16'hFFDB;
        rom[32][94] = 16'hFFFE;
        rom[32][95] = 16'h0003;
        rom[32][96] = 16'hFFC8;
        rom[32][97] = 16'h0023;
        rom[32][98] = 16'h001C;
        rom[32][99] = 16'h0015;
        rom[32][100] = 16'hFFD5;
        rom[32][101] = 16'hFFF8;
        rom[32][102] = 16'h0007;
        rom[32][103] = 16'h000B;
        rom[32][104] = 16'hFFF6;
        rom[32][105] = 16'h000B;
        rom[32][106] = 16'h002E;
        rom[32][107] = 16'hFFCA;
        rom[32][108] = 16'hFFEE;
        rom[32][109] = 16'h0009;
        rom[32][110] = 16'h001B;
        rom[32][111] = 16'hFFE0;
        rom[32][112] = 16'hFFCD;
        rom[32][113] = 16'hFFD4;
        rom[32][114] = 16'h0035;
        rom[32][115] = 16'hFFD7;
        rom[32][116] = 16'h0007;
        rom[32][117] = 16'h0019;
        rom[32][118] = 16'hFFF7;
        rom[32][119] = 16'h0008;
        rom[32][120] = 16'hFFEA;
        rom[32][121] = 16'hFFF6;
        rom[32][122] = 16'h000E;
        rom[32][123] = 16'h0024;
        rom[32][124] = 16'h0007;
        rom[32][125] = 16'hFFEF;
        rom[32][126] = 16'hFFF8;
        rom[32][127] = 16'hFFE2;
        rom[33][0] = 16'hFFC6;
        rom[33][1] = 16'hFFD7;
        rom[33][2] = 16'h0011;
        rom[33][3] = 16'h001B;
        rom[33][4] = 16'hFFE8;
        rom[33][5] = 16'hFFC6;
        rom[33][6] = 16'hFFE4;
        rom[33][7] = 16'h0016;
        rom[33][8] = 16'hFFB2;
        rom[33][9] = 16'h0005;
        rom[33][10] = 16'h001B;
        rom[33][11] = 16'hFFEA;
        rom[33][12] = 16'hFFC7;
        rom[33][13] = 16'h0014;
        rom[33][14] = 16'hFFD8;
        rom[33][15] = 16'hFFF2;
        rom[33][16] = 16'hFFD3;
        rom[33][17] = 16'h0012;
        rom[33][18] = 16'hFFE5;
        rom[33][19] = 16'h0039;
        rom[33][20] = 16'h0007;
        rom[33][21] = 16'h001C;
        rom[33][22] = 16'h001F;
        rom[33][23] = 16'hFFEE;
        rom[33][24] = 16'h0007;
        rom[33][25] = 16'hFFDA;
        rom[33][26] = 16'h001C;
        rom[33][27] = 16'h0003;
        rom[33][28] = 16'h000C;
        rom[33][29] = 16'h0007;
        rom[33][30] = 16'h0007;
        rom[33][31] = 16'h0019;
        rom[33][32] = 16'h0029;
        rom[33][33] = 16'h0002;
        rom[33][34] = 16'hFFFD;
        rom[33][35] = 16'hFFF6;
        rom[33][36] = 16'hFFEC;
        rom[33][37] = 16'h000A;
        rom[33][38] = 16'h000A;
        rom[33][39] = 16'hFFEC;
        rom[33][40] = 16'h0015;
        rom[33][41] = 16'hFFE2;
        rom[33][42] = 16'hFFE2;
        rom[33][43] = 16'hFFEA;
        rom[33][44] = 16'h0001;
        rom[33][45] = 16'hFFF8;
        rom[33][46] = 16'hFFE0;
        rom[33][47] = 16'hFFC8;
        rom[33][48] = 16'hFFE4;
        rom[33][49] = 16'hFFB0;
        rom[33][50] = 16'hFFF4;
        rom[33][51] = 16'h0006;
        rom[33][52] = 16'h0010;
        rom[33][53] = 16'hFFD3;
        rom[33][54] = 16'h001B;
        rom[33][55] = 16'hFFE5;
        rom[33][56] = 16'h001A;
        rom[33][57] = 16'hFFEE;
        rom[33][58] = 16'h0004;
        rom[33][59] = 16'hFFFA;
        rom[33][60] = 16'hFFEA;
        rom[33][61] = 16'h0014;
        rom[33][62] = 16'hFFC8;
        rom[33][63] = 16'hFFF7;
        rom[33][64] = 16'h0034;
        rom[33][65] = 16'hFFFD;
        rom[33][66] = 16'hFFFE;
        rom[33][67] = 16'hFFE5;
        rom[33][68] = 16'hFFDD;
        rom[33][69] = 16'hFFD0;
        rom[33][70] = 16'hFFE0;
        rom[33][71] = 16'hFFFC;
        rom[33][72] = 16'hFFEA;
        rom[33][73] = 16'hFFF9;
        rom[33][74] = 16'hFFF9;
        rom[33][75] = 16'h0016;
        rom[33][76] = 16'hFFF9;
        rom[33][77] = 16'h0012;
        rom[33][78] = 16'hFFE0;
        rom[33][79] = 16'hFFBF;
        rom[33][80] = 16'hFFF9;
        rom[33][81] = 16'hFFE1;
        rom[33][82] = 16'h0007;
        rom[33][83] = 16'h0015;
        rom[33][84] = 16'hFFA3;
        rom[33][85] = 16'h0014;
        rom[33][86] = 16'h0016;
        rom[33][87] = 16'h0014;
        rom[33][88] = 16'h0026;
        rom[33][89] = 16'h0009;
        rom[33][90] = 16'h0011;
        rom[33][91] = 16'hFFEF;
        rom[33][92] = 16'hFFEA;
        rom[33][93] = 16'hFFEC;
        rom[33][94] = 16'h0020;
        rom[33][95] = 16'hFFD2;
        rom[33][96] = 16'hFFC4;
        rom[33][97] = 16'hFFF8;
        rom[33][98] = 16'h0032;
        rom[33][99] = 16'hFFD5;
        rom[33][100] = 16'h0002;
        rom[33][101] = 16'h0005;
        rom[33][102] = 16'hFFE0;
        rom[33][103] = 16'hFFC8;
        rom[33][104] = 16'h0020;
        rom[33][105] = 16'h0003;
        rom[33][106] = 16'h0021;
        rom[33][107] = 16'hFF9E;
        rom[33][108] = 16'hFFFE;
        rom[33][109] = 16'h0003;
        rom[33][110] = 16'h0007;
        rom[33][111] = 16'hFFE5;
        rom[33][112] = 16'hFFF7;
        rom[33][113] = 16'h0000;
        rom[33][114] = 16'hFFF8;
        rom[33][115] = 16'hFFF9;
        rom[33][116] = 16'hFFF4;
        rom[33][117] = 16'hFFDC;
        rom[33][118] = 16'hFFF2;
        rom[33][119] = 16'h0001;
        rom[33][120] = 16'hFFEF;
        rom[33][121] = 16'hFFFD;
        rom[33][122] = 16'hFFC8;
        rom[33][123] = 16'hFFF7;
        rom[33][124] = 16'h000D;
        rom[33][125] = 16'hFFEB;
        rom[33][126] = 16'hFFE3;
        rom[33][127] = 16'hFFDA;
        rom[34][0] = 16'h002C;
        rom[34][1] = 16'hFFEA;
        rom[34][2] = 16'hFFD3;
        rom[34][3] = 16'h0007;
        rom[34][4] = 16'hFFFB;
        rom[34][5] = 16'hFFEE;
        rom[34][6] = 16'h000A;
        rom[34][7] = 16'h0002;
        rom[34][8] = 16'h0002;
        rom[34][9] = 16'h0016;
        rom[34][10] = 16'h0007;
        rom[34][11] = 16'h000B;
        rom[34][12] = 16'h0017;
        rom[34][13] = 16'h0004;
        rom[34][14] = 16'h0016;
        rom[34][15] = 16'hFFF4;
        rom[34][16] = 16'hFFD0;
        rom[34][17] = 16'hFFD7;
        rom[34][18] = 16'h001E;
        rom[34][19] = 16'hFFE0;
        rom[34][20] = 16'hFFF4;
        rom[34][21] = 16'h0010;
        rom[34][22] = 16'hFFD8;
        rom[34][23] = 16'h0018;
        rom[34][24] = 16'h0007;
        rom[34][25] = 16'hFFE7;
        rom[34][26] = 16'hFFDD;
        rom[34][27] = 16'hFFEA;
        rom[34][28] = 16'hFFE4;
        rom[34][29] = 16'hFFC1;
        rom[34][30] = 16'h0006;
        rom[34][31] = 16'hFFD9;
        rom[34][32] = 16'hFFAF;
        rom[34][33] = 16'h000E;
        rom[34][34] = 16'h0010;
        rom[34][35] = 16'hFFF3;
        rom[34][36] = 16'h0007;
        rom[34][37] = 16'hFFF4;
        rom[34][38] = 16'h000D;
        rom[34][39] = 16'hFFDC;
        rom[34][40] = 16'hFFC3;
        rom[34][41] = 16'h0016;
        rom[34][42] = 16'h0000;
        rom[34][43] = 16'h003D;
        rom[34][44] = 16'hFFE1;
        rom[34][45] = 16'hFFE5;
        rom[34][46] = 16'hFFFB;
        rom[34][47] = 16'hFFF8;
        rom[34][48] = 16'hFFE8;
        rom[34][49] = 16'h0001;
        rom[34][50] = 16'hFFE5;
        rom[34][51] = 16'h0005;
        rom[34][52] = 16'h0004;
        rom[34][53] = 16'hFFF1;
        rom[34][54] = 16'hFFB6;
        rom[34][55] = 16'hFFFA;
        rom[34][56] = 16'hFFDC;
        rom[34][57] = 16'hFFE3;
        rom[34][58] = 16'h001C;
        rom[34][59] = 16'h000D;
        rom[34][60] = 16'hFFF6;
        rom[34][61] = 16'hFFD3;
        rom[34][62] = 16'hFFDF;
        rom[34][63] = 16'h0022;
        rom[34][64] = 16'hFFDE;
        rom[34][65] = 16'h0011;
        rom[34][66] = 16'hFFFE;
        rom[34][67] = 16'hFFFB;
        rom[34][68] = 16'h0005;
        rom[34][69] = 16'h0013;
        rom[34][70] = 16'hFFE1;
        rom[34][71] = 16'h001A;
        rom[34][72] = 16'hFFF8;
        rom[34][73] = 16'hFFDC;
        rom[34][74] = 16'h0022;
        rom[34][75] = 16'h0032;
        rom[34][76] = 16'h002C;
        rom[34][77] = 16'h0011;
        rom[34][78] = 16'hFF9F;
        rom[34][79] = 16'h0016;
        rom[34][80] = 16'hFFFF;
        rom[34][81] = 16'h0002;
        rom[34][82] = 16'h0002;
        rom[34][83] = 16'hFFD1;
        rom[34][84] = 16'h0009;
        rom[34][85] = 16'hFFDA;
        rom[34][86] = 16'hFFCC;
        rom[34][87] = 16'h0026;
        rom[34][88] = 16'hFFD0;
        rom[34][89] = 16'hFFC1;
        rom[34][90] = 16'hFFCD;
        rom[34][91] = 16'h0004;
        rom[34][92] = 16'h002C;
        rom[34][93] = 16'h000C;
        rom[34][94] = 16'hFFFC;
        rom[34][95] = 16'h0004;
        rom[34][96] = 16'h001D;
        rom[34][97] = 16'hFFF9;
        rom[34][98] = 16'hFFFB;
        rom[34][99] = 16'hFFFD;
        rom[34][100] = 16'hFFD5;
        rom[34][101] = 16'hFFEE;
        rom[34][102] = 16'h001F;
        rom[34][103] = 16'h0027;
        rom[34][104] = 16'h0000;
        rom[34][105] = 16'hFFE1;
        rom[34][106] = 16'hFFDE;
        rom[34][107] = 16'h0008;
        rom[34][108] = 16'hFFE1;
        rom[34][109] = 16'h0015;
        rom[34][110] = 16'hFFE6;
        rom[34][111] = 16'hFFF1;
        rom[34][112] = 16'h0025;
        rom[34][113] = 16'h0011;
        rom[34][114] = 16'h0025;
        rom[34][115] = 16'h0002;
        rom[34][116] = 16'h0022;
        rom[34][117] = 16'h0006;
        rom[34][118] = 16'hFFEA;
        rom[34][119] = 16'hFFE4;
        rom[34][120] = 16'h0006;
        rom[34][121] = 16'h0010;
        rom[34][122] = 16'h003C;
        rom[34][123] = 16'h001B;
        rom[34][124] = 16'hFFF0;
        rom[34][125] = 16'h002E;
        rom[34][126] = 16'h002E;
        rom[34][127] = 16'h0029;
        rom[35][0] = 16'h0006;
        rom[35][1] = 16'hFFF2;
        rom[35][2] = 16'h0007;
        rom[35][3] = 16'hFFF9;
        rom[35][4] = 16'h000D;
        rom[35][5] = 16'hFFBC;
        rom[35][6] = 16'h0003;
        rom[35][7] = 16'hFFCD;
        rom[35][8] = 16'hFFFE;
        rom[35][9] = 16'h000C;
        rom[35][10] = 16'hFFEB;
        rom[35][11] = 16'h000A;
        rom[35][12] = 16'h0007;
        rom[35][13] = 16'h0007;
        rom[35][14] = 16'hFFED;
        rom[35][15] = 16'h002E;
        rom[35][16] = 16'hFFEA;
        rom[35][17] = 16'hFFC3;
        rom[35][18] = 16'hFFFF;
        rom[35][19] = 16'hFFE9;
        rom[35][20] = 16'hFFF4;
        rom[35][21] = 16'hFFF2;
        rom[35][22] = 16'h0004;
        rom[35][23] = 16'hFFDC;
        rom[35][24] = 16'hFFF0;
        rom[35][25] = 16'hFFD2;
        rom[35][26] = 16'hFFEF;
        rom[35][27] = 16'h0003;
        rom[35][28] = 16'hFFEB;
        rom[35][29] = 16'h000C;
        rom[35][30] = 16'h000A;
        rom[35][31] = 16'hFFF6;
        rom[35][32] = 16'h0002;
        rom[35][33] = 16'h0004;
        rom[35][34] = 16'h000D;
        rom[35][35] = 16'hFFF6;
        rom[35][36] = 16'hFFF6;
        rom[35][37] = 16'h001B;
        rom[35][38] = 16'h0007;
        rom[35][39] = 16'hFFF0;
        rom[35][40] = 16'h0000;
        rom[35][41] = 16'h000E;
        rom[35][42] = 16'hFFFC;
        rom[35][43] = 16'hFFEE;
        rom[35][44] = 16'h0019;
        rom[35][45] = 16'hFFE5;
        rom[35][46] = 16'h001A;
        rom[35][47] = 16'hFFA5;
        rom[35][48] = 16'h000B;
        rom[35][49] = 16'hFFC3;
        rom[35][50] = 16'hFFFC;
        rom[35][51] = 16'hFFEA;
        rom[35][52] = 16'h0002;
        rom[35][53] = 16'hFFEC;
        rom[35][54] = 16'hFFEF;
        rom[35][55] = 16'hFFFF;
        rom[35][56] = 16'hFFE5;
        rom[35][57] = 16'hFFEC;
        rom[35][58] = 16'hFFFE;
        rom[35][59] = 16'h0008;
        rom[35][60] = 16'h0005;
        rom[35][61] = 16'hFFEB;
        rom[35][62] = 16'hFFD6;
        rom[35][63] = 16'hFFA4;
        rom[35][64] = 16'h000E;
        rom[35][65] = 16'h0000;
        rom[35][66] = 16'hFFF8;
        rom[35][67] = 16'hFFDC;
        rom[35][68] = 16'hFFE2;
        rom[35][69] = 16'hFFDC;
        rom[35][70] = 16'h0005;
        rom[35][71] = 16'h0001;
        rom[35][72] = 16'h0015;
        rom[35][73] = 16'h0009;
        rom[35][74] = 16'hFFC3;
        rom[35][75] = 16'hFFFD;
        rom[35][76] = 16'hFFF9;
        rom[35][77] = 16'h0009;
        rom[35][78] = 16'hFFFC;
        rom[35][79] = 16'h0033;
        rom[35][80] = 16'hFFA9;
        rom[35][81] = 16'h0016;
        rom[35][82] = 16'hFFC5;
        rom[35][83] = 16'h0038;
        rom[35][84] = 16'h000B;
        rom[35][85] = 16'h0002;
        rom[35][86] = 16'h0002;
        rom[35][87] = 16'h000C;
        rom[35][88] = 16'hFFF8;
        rom[35][89] = 16'h001B;
        rom[35][90] = 16'hFFCD;
        rom[35][91] = 16'hFFED;
        rom[35][92] = 16'h0018;
        rom[35][93] = 16'hFFCB;
        rom[35][94] = 16'hFFCB;
        rom[35][95] = 16'hFFB5;
        rom[35][96] = 16'hFFC0;
        rom[35][97] = 16'h000D;
        rom[35][98] = 16'hFFA6;
        rom[35][99] = 16'h000F;
        rom[35][100] = 16'hFFD7;
        rom[35][101] = 16'hFFE4;
        rom[35][102] = 16'hFFEF;
        rom[35][103] = 16'hFFF0;
        rom[35][104] = 16'h0002;
        rom[35][105] = 16'hFFFF;
        rom[35][106] = 16'h0016;
        rom[35][107] = 16'h0022;
        rom[35][108] = 16'hFFF4;
        rom[35][109] = 16'hFFF8;
        rom[35][110] = 16'h000B;
        rom[35][111] = 16'hFFC7;
        rom[35][112] = 16'hFFCD;
        rom[35][113] = 16'h000B;
        rom[35][114] = 16'hFFE6;
        rom[35][115] = 16'hFFE1;
        rom[35][116] = 16'h0012;
        rom[35][117] = 16'hFFEE;
        rom[35][118] = 16'hFFDA;
        rom[35][119] = 16'h0018;
        rom[35][120] = 16'h0016;
        rom[35][121] = 16'hFFDE;
        rom[35][122] = 16'h000D;
        rom[35][123] = 16'h002B;
        rom[35][124] = 16'h0011;
        rom[35][125] = 16'h0011;
        rom[35][126] = 16'hFFEF;
        rom[35][127] = 16'hFFFE;
        rom[36][0] = 16'h0037;
        rom[36][1] = 16'hFFD7;
        rom[36][2] = 16'h0002;
        rom[36][3] = 16'hFFF5;
        rom[36][4] = 16'h0002;
        rom[36][5] = 16'hFFF5;
        rom[36][6] = 16'hFFEE;
        rom[36][7] = 16'h0007;
        rom[36][8] = 16'h001A;
        rom[36][9] = 16'hFFE2;
        rom[36][10] = 16'h0020;
        rom[36][11] = 16'h001B;
        rom[36][12] = 16'h0016;
        rom[36][13] = 16'h0021;
        rom[36][14] = 16'hFFE9;
        rom[36][15] = 16'hFFDE;
        rom[36][16] = 16'h000F;
        rom[36][17] = 16'hFFD9;
        rom[36][18] = 16'h000F;
        rom[36][19] = 16'hFFDC;
        rom[36][20] = 16'hFFF9;
        rom[36][21] = 16'hFFF5;
        rom[36][22] = 16'hFFC7;
        rom[36][23] = 16'h0017;
        rom[36][24] = 16'hFFF2;
        rom[36][25] = 16'h005C;
        rom[36][26] = 16'h0007;
        rom[36][27] = 16'hFFE9;
        rom[36][28] = 16'hFFCD;
        rom[36][29] = 16'hFFC1;
        rom[36][30] = 16'h005A;
        rom[36][31] = 16'h0049;
        rom[36][32] = 16'h0011;
        rom[36][33] = 16'hFFE4;
        rom[36][34] = 16'hFFF9;
        rom[36][35] = 16'hFFE1;
        rom[36][36] = 16'h001B;
        rom[36][37] = 16'hFFC3;
        rom[36][38] = 16'hFFEF;
        rom[36][39] = 16'hFFFE;
        rom[36][40] = 16'h0007;
        rom[36][41] = 16'h0013;
        rom[36][42] = 16'h0018;
        rom[36][43] = 16'hFFC2;
        rom[36][44] = 16'h001F;
        rom[36][45] = 16'hFFE5;
        rom[36][46] = 16'h0014;
        rom[36][47] = 16'hFFCF;
        rom[36][48] = 16'h0014;
        rom[36][49] = 16'h001B;
        rom[36][50] = 16'hFFEA;
        rom[36][51] = 16'h0020;
        rom[36][52] = 16'hFFB3;
        rom[36][53] = 16'hFFEE;
        rom[36][54] = 16'hFFD8;
        rom[36][55] = 16'h0009;
        rom[36][56] = 16'h0011;
        rom[36][57] = 16'hFFE1;
        rom[36][58] = 16'hFFDB;
        rom[36][59] = 16'h0011;
        rom[36][60] = 16'h0003;
        rom[36][61] = 16'h0033;
        rom[36][62] = 16'hFFE8;
        rom[36][63] = 16'hFFDC;
        rom[36][64] = 16'hFFF0;
        rom[36][65] = 16'h0008;
        rom[36][66] = 16'hFFCA;
        rom[36][67] = 16'h000A;
        rom[36][68] = 16'h0006;
        rom[36][69] = 16'hFFE9;
        rom[36][70] = 16'hFFFC;
        rom[36][71] = 16'hFF9D;
        rom[36][72] = 16'h0007;
        rom[36][73] = 16'h0013;
        rom[36][74] = 16'h0034;
        rom[36][75] = 16'hFFCF;
        rom[36][76] = 16'h000B;
        rom[36][77] = 16'h002F;
        rom[36][78] = 16'hFFFD;
        rom[36][79] = 16'h000E;
        rom[36][80] = 16'hFFD1;
        rom[36][81] = 16'hFFDF;
        rom[36][82] = 16'hFFEE;
        rom[36][83] = 16'h0015;
        rom[36][84] = 16'hFFFC;
        rom[36][85] = 16'hFFC0;
        rom[36][86] = 16'h002A;
        rom[36][87] = 16'hFFD0;
        rom[36][88] = 16'h001B;
        rom[36][89] = 16'hFFBE;
        rom[36][90] = 16'h001C;
        rom[36][91] = 16'hFFF5;
        rom[36][92] = 16'hFFFE;
        rom[36][93] = 16'hFFCA;
        rom[36][94] = 16'hFFD6;
        rom[36][95] = 16'h0002;
        rom[36][96] = 16'hFFB5;
        rom[36][97] = 16'h001C;
        rom[36][98] = 16'h0016;
        rom[36][99] = 16'h0003;
        rom[36][100] = 16'hFFD7;
        rom[36][101] = 16'hFFDA;
        rom[36][102] = 16'hFFFB;
        rom[36][103] = 16'hFFFD;
        rom[36][104] = 16'h004B;
        rom[36][105] = 16'h0041;
        rom[36][106] = 16'hFFCE;
        rom[36][107] = 16'h0007;
        rom[36][108] = 16'hFFF4;
        rom[36][109] = 16'hFFE7;
        rom[36][110] = 16'h0003;
        rom[36][111] = 16'hFFDB;
        rom[36][112] = 16'hFFEF;
        rom[36][113] = 16'h0029;
        rom[36][114] = 16'h0021;
        rom[36][115] = 16'h001D;
        rom[36][116] = 16'hFFE9;
        rom[36][117] = 16'hFFC8;
        rom[36][118] = 16'hFFF1;
        rom[36][119] = 16'hFFEF;
        rom[36][120] = 16'h004A;
        rom[36][121] = 16'hFFEE;
        rom[36][122] = 16'hFFFC;
        rom[36][123] = 16'hFFF8;
        rom[36][124] = 16'hFFCE;
        rom[36][125] = 16'h0038;
        rom[36][126] = 16'hFFE5;
        rom[36][127] = 16'hFFE5;
        rom[37][0] = 16'h0002;
        rom[37][1] = 16'hFFF0;
        rom[37][2] = 16'hFFD0;
        rom[37][3] = 16'hFFF9;
        rom[37][4] = 16'hFFF9;
        rom[37][5] = 16'hFFE2;
        rom[37][6] = 16'hFFE5;
        rom[37][7] = 16'h0037;
        rom[37][8] = 16'hFFE0;
        rom[37][9] = 16'hFFEB;
        rom[37][10] = 16'h0017;
        rom[37][11] = 16'hFFEF;
        rom[37][12] = 16'h000C;
        rom[37][13] = 16'h0011;
        rom[37][14] = 16'hFFD7;
        rom[37][15] = 16'hFFCE;
        rom[37][16] = 16'h001B;
        rom[37][17] = 16'h0037;
        rom[37][18] = 16'h0016;
        rom[37][19] = 16'h0040;
        rom[37][20] = 16'h0020;
        rom[37][21] = 16'hFFFB;
        rom[37][22] = 16'h0011;
        rom[37][23] = 16'h001A;
        rom[37][24] = 16'hFFBA;
        rom[37][25] = 16'hFFAC;
        rom[37][26] = 16'hFFEF;
        rom[37][27] = 16'hFFFE;
        rom[37][28] = 16'h0013;
        rom[37][29] = 16'h0016;
        rom[37][30] = 16'h0011;
        rom[37][31] = 16'hFFD8;
        rom[37][32] = 16'hFFE9;
        rom[37][33] = 16'h0035;
        rom[37][34] = 16'hFFC7;
        rom[37][35] = 16'hFFFE;
        rom[37][36] = 16'h000E;
        rom[37][37] = 16'hFFE6;
        rom[37][38] = 16'h0024;
        rom[37][39] = 16'h003E;
        rom[37][40] = 16'hFFF5;
        rom[37][41] = 16'h0003;
        rom[37][42] = 16'hFFF4;
        rom[37][43] = 16'hFFFE;
        rom[37][44] = 16'h0029;
        rom[37][45] = 16'h0007;
        rom[37][46] = 16'h000D;
        rom[37][47] = 16'hFFCF;
        rom[37][48] = 16'hFFDA;
        rom[37][49] = 16'hFFDE;
        rom[37][50] = 16'hFFC0;
        rom[37][51] = 16'h0015;
        rom[37][52] = 16'hFFF6;
        rom[37][53] = 16'hFFF4;
        rom[37][54] = 16'h000B;
        rom[37][55] = 16'hFFEF;
        rom[37][56] = 16'hFFFD;
        rom[37][57] = 16'h0016;
        rom[37][58] = 16'h0009;
        rom[37][59] = 16'h0018;
        rom[37][60] = 16'h0033;
        rom[37][61] = 16'h000C;
        rom[37][62] = 16'h0008;
        rom[37][63] = 16'hFFCB;
        rom[37][64] = 16'hFFD7;
        rom[37][65] = 16'h0034;
        rom[37][66] = 16'hFFD6;
        rom[37][67] = 16'hFFEF;
        rom[37][68] = 16'hFFFB;
        rom[37][69] = 16'hFFEF;
        rom[37][70] = 16'hFFB8;
        rom[37][71] = 16'hFFF3;
        rom[37][72] = 16'hFFF9;
        rom[37][73] = 16'hFFE4;
        rom[37][74] = 16'hFFEB;
        rom[37][75] = 16'h0005;
        rom[37][76] = 16'hFFB8;
        rom[37][77] = 16'h0034;
        rom[37][78] = 16'h0005;
        rom[37][79] = 16'h0029;
        rom[37][80] = 16'hFFB5;
        rom[37][81] = 16'h000C;
        rom[37][82] = 16'hFFEC;
        rom[37][83] = 16'h000E;
        rom[37][84] = 16'h0001;
        rom[37][85] = 16'hFFFC;
        rom[37][86] = 16'hFFF6;
        rom[37][87] = 16'hFFEF;
        rom[37][88] = 16'h0002;
        rom[37][89] = 16'h000E;
        rom[37][90] = 16'h000F;
        rom[37][91] = 16'h0001;
        rom[37][92] = 16'h0062;
        rom[37][93] = 16'h0021;
        rom[37][94] = 16'h003B;
        rom[37][95] = 16'h0009;
        rom[37][96] = 16'h0011;
        rom[37][97] = 16'h0014;
        rom[37][98] = 16'h001B;
        rom[37][99] = 16'h0038;
        rom[37][100] = 16'hFFF8;
        rom[37][101] = 16'h0018;
        rom[37][102] = 16'hFFBA;
        rom[37][103] = 16'hFFF4;
        rom[37][104] = 16'hFFDD;
        rom[37][105] = 16'hFFEE;
        rom[37][106] = 16'hFFE1;
        rom[37][107] = 16'hFFED;
        rom[37][108] = 16'h0005;
        rom[37][109] = 16'h0006;
        rom[37][110] = 16'hFFEF;
        rom[37][111] = 16'h0018;
        rom[37][112] = 16'h0038;
        rom[37][113] = 16'hFFFE;
        rom[37][114] = 16'h0016;
        rom[37][115] = 16'h003A;
        rom[37][116] = 16'hFFFE;
        rom[37][117] = 16'h0037;
        rom[37][118] = 16'hFFC6;
        rom[37][119] = 16'h0009;
        rom[37][120] = 16'hFFC7;
        rom[37][121] = 16'h0011;
        rom[37][122] = 16'hFFF6;
        rom[37][123] = 16'hFFB0;
        rom[37][124] = 16'h001B;
        rom[37][125] = 16'hFFF6;
        rom[37][126] = 16'hFFFB;
        rom[37][127] = 16'h000F;
        rom[38][0] = 16'hFFF0;
        rom[38][1] = 16'hFFFF;
        rom[38][2] = 16'hFFF6;
        rom[38][3] = 16'hFFE5;
        rom[38][4] = 16'hFFF9;
        rom[38][5] = 16'hFFB2;
        rom[38][6] = 16'hFFE1;
        rom[38][7] = 16'h0016;
        rom[38][8] = 16'hFFF7;
        rom[38][9] = 16'hFFD2;
        rom[38][10] = 16'hFFE5;
        rom[38][11] = 16'hFFF2;
        rom[38][12] = 16'h0012;
        rom[38][13] = 16'h0011;
        rom[38][14] = 16'hFFDA;
        rom[38][15] = 16'h0003;
        rom[38][16] = 16'hFFB1;
        rom[38][17] = 16'h0027;
        rom[38][18] = 16'h001A;
        rom[38][19] = 16'hFFE5;
        rom[38][20] = 16'h0015;
        rom[38][21] = 16'h0012;
        rom[38][22] = 16'h0036;
        rom[38][23] = 16'h001E;
        rom[38][24] = 16'h0015;
        rom[38][25] = 16'hFFC8;
        rom[38][26] = 16'h0011;
        rom[38][27] = 16'hFFB4;
        rom[38][28] = 16'hFFD8;
        rom[38][29] = 16'h0012;
        rom[38][30] = 16'hFFE4;
        rom[38][31] = 16'hFFFC;
        rom[38][32] = 16'h0011;
        rom[38][33] = 16'h0003;
        rom[38][34] = 16'hFFEC;
        rom[38][35] = 16'h000D;
        rom[38][36] = 16'hFFFB;
        rom[38][37] = 16'h0046;
        rom[38][38] = 16'h001B;
        rom[38][39] = 16'hFFF6;
        rom[38][40] = 16'hFFE9;
        rom[38][41] = 16'hFFFF;
        rom[38][42] = 16'h003C;
        rom[38][43] = 16'hFFD3;
        rom[38][44] = 16'h0033;
        rom[38][45] = 16'h000D;
        rom[38][46] = 16'h0016;
        rom[38][47] = 16'hFFE6;
        rom[38][48] = 16'h000C;
        rom[38][49] = 16'hFFD5;
        rom[38][50] = 16'h0024;
        rom[38][51] = 16'hFFEF;
        rom[38][52] = 16'hFFE1;
        rom[38][53] = 16'hFFE1;
        rom[38][54] = 16'hFFE5;
        rom[38][55] = 16'hFFE0;
        rom[38][56] = 16'h0002;
        rom[38][57] = 16'hFFE4;
        rom[38][58] = 16'h0018;
        rom[38][59] = 16'hFFED;
        rom[38][60] = 16'hFFBD;
        rom[38][61] = 16'hFFDC;
        rom[38][62] = 16'h0003;
        rom[38][63] = 16'hFFD7;
        rom[38][64] = 16'hFFE3;
        rom[38][65] = 16'hFFFD;
        rom[38][66] = 16'h0001;
        rom[38][67] = 16'hFFCC;
        rom[38][68] = 16'hFFF9;
        rom[38][69] = 16'hFFD2;
        rom[38][70] = 16'h001C;
        rom[38][71] = 16'hFFB5;
        rom[38][72] = 16'hFFFE;
        rom[38][73] = 16'hFFF9;
        rom[38][74] = 16'h001F;
        rom[38][75] = 16'hFFF9;
        rom[38][76] = 16'hFFF0;
        rom[38][77] = 16'hFFFE;
        rom[38][78] = 16'hFFF9;
        rom[38][79] = 16'hFFEF;
        rom[38][80] = 16'hFFF3;
        rom[38][81] = 16'h0041;
        rom[38][82] = 16'hFFD3;
        rom[38][83] = 16'h000C;
        rom[38][84] = 16'h0010;
        rom[38][85] = 16'hFFC0;
        rom[38][86] = 16'hFFDB;
        rom[38][87] = 16'hFFE3;
        rom[38][88] = 16'hFFDE;
        rom[38][89] = 16'h0007;
        rom[38][90] = 16'hFFE4;
        rom[38][91] = 16'hFFEA;
        rom[38][92] = 16'h0044;
        rom[38][93] = 16'h0041;
        rom[38][94] = 16'h000B;
        rom[38][95] = 16'h0040;
        rom[38][96] = 16'hFFF7;
        rom[38][97] = 16'hFFF6;
        rom[38][98] = 16'hFFAE;
        rom[38][99] = 16'h0020;
        rom[38][100] = 16'hFFF4;
        rom[38][101] = 16'hFFFC;
        rom[38][102] = 16'hFFF5;
        rom[38][103] = 16'h0007;
        rom[38][104] = 16'hFFE1;
        rom[38][105] = 16'hFFFE;
        rom[38][106] = 16'hFFE1;
        rom[38][107] = 16'h0016;
        rom[38][108] = 16'hFFC9;
        rom[38][109] = 16'h002E;
        rom[38][110] = 16'hFFD9;
        rom[38][111] = 16'hFFDC;
        rom[38][112] = 16'hFFF6;
        rom[38][113] = 16'hFFE7;
        rom[38][114] = 16'h000B;
        rom[38][115] = 16'hFFEA;
        rom[38][116] = 16'h0001;
        rom[38][117] = 16'h0002;
        rom[38][118] = 16'hFFCA;
        rom[38][119] = 16'h0029;
        rom[38][120] = 16'hFFE5;
        rom[38][121] = 16'hFFC3;
        rom[38][122] = 16'hFFF0;
        rom[38][123] = 16'h0021;
        rom[38][124] = 16'h0011;
        rom[38][125] = 16'hFFF8;
        rom[38][126] = 16'h0009;
        rom[38][127] = 16'hFFF1;
        rom[39][0] = 16'hFFCE;
        rom[39][1] = 16'h000E;
        rom[39][2] = 16'h0021;
        rom[39][3] = 16'hFFE6;
        rom[39][4] = 16'h0007;
        rom[39][5] = 16'h001D;
        rom[39][6] = 16'h0015;
        rom[39][7] = 16'h001F;
        rom[39][8] = 16'hFFFC;
        rom[39][9] = 16'hFFE2;
        rom[39][10] = 16'hFFD3;
        rom[39][11] = 16'h0002;
        rom[39][12] = 16'hFFE7;
        rom[39][13] = 16'hFFEA;
        rom[39][14] = 16'h0021;
        rom[39][15] = 16'hFFF0;
        rom[39][16] = 16'h0003;
        rom[39][17] = 16'hFFF1;
        rom[39][18] = 16'hFFFF;
        rom[39][19] = 16'hFFE7;
        rom[39][20] = 16'h0014;
        rom[39][21] = 16'h0016;
        rom[39][22] = 16'hFFC6;
        rom[39][23] = 16'hFFB0;
        rom[39][24] = 16'hFFE3;
        rom[39][25] = 16'h001F;
        rom[39][26] = 16'hFFF4;
        rom[39][27] = 16'hFFF6;
        rom[39][28] = 16'hFFEF;
        rom[39][29] = 16'hFFE9;
        rom[39][30] = 16'h000C;
        rom[39][31] = 16'hFFF3;
        rom[39][32] = 16'hFFC3;
        rom[39][33] = 16'hFFE0;
        rom[39][34] = 16'h000D;
        rom[39][35] = 16'hFFDA;
        rom[39][36] = 16'h0005;
        rom[39][37] = 16'h0030;
        rom[39][38] = 16'h000E;
        rom[39][39] = 16'hFFFE;
        rom[39][40] = 16'hFFF6;
        rom[39][41] = 16'h0012;
        rom[39][42] = 16'hFFEE;
        rom[39][43] = 16'hFFFF;
        rom[39][44] = 16'hFFDB;
        rom[39][45] = 16'hFFDE;
        rom[39][46] = 16'h0019;
        rom[39][47] = 16'hFFF4;
        rom[39][48] = 16'hFFD2;
        rom[39][49] = 16'hFFF9;
        rom[39][50] = 16'h000B;
        rom[39][51] = 16'hFFF3;
        rom[39][52] = 16'h001A;
        rom[39][53] = 16'h000C;
        rom[39][54] = 16'hFFEA;
        rom[39][55] = 16'h0017;
        rom[39][56] = 16'hFFDC;
        rom[39][57] = 16'hFFB5;
        rom[39][58] = 16'h0017;
        rom[39][59] = 16'hFFE5;
        rom[39][60] = 16'h001D;
        rom[39][61] = 16'hFFE9;
        rom[39][62] = 16'hFFF3;
        rom[39][63] = 16'h0017;
        rom[39][64] = 16'h000E;
        rom[39][65] = 16'h0016;
        rom[39][66] = 16'h001D;
        rom[39][67] = 16'h000A;
        rom[39][68] = 16'h0013;
        rom[39][69] = 16'h0033;
        rom[39][70] = 16'h0016;
        rom[39][71] = 16'h001E;
        rom[39][72] = 16'hFFC6;
        rom[39][73] = 16'h000E;
        rom[39][74] = 16'h0013;
        rom[39][75] = 16'h001B;
        rom[39][76] = 16'h0000;
        rom[39][77] = 16'h0016;
        rom[39][78] = 16'hFFEB;
        rom[39][79] = 16'h002E;
        rom[39][80] = 16'h002A;
        rom[39][81] = 16'hFFFA;
        rom[39][82] = 16'h001F;
        rom[39][83] = 16'hFFFC;
        rom[39][84] = 16'hFFF4;
        rom[39][85] = 16'h0016;
        rom[39][86] = 16'hFFEC;
        rom[39][87] = 16'h0016;
        rom[39][88] = 16'hFFE1;
        rom[39][89] = 16'h000A;
        rom[39][90] = 16'h0002;
        rom[39][91] = 16'hFFF0;
        rom[39][92] = 16'h0041;
        rom[39][93] = 16'hFFC3;
        rom[39][94] = 16'h0024;
        rom[39][95] = 16'hFFEA;
        rom[39][96] = 16'hFFE5;
        rom[39][97] = 16'hFFE0;
        rom[39][98] = 16'hFFDC;
        rom[39][99] = 16'h0009;
        rom[39][100] = 16'hFFAB;
        rom[39][101] = 16'hFFE1;
        rom[39][102] = 16'hFFFE;
        rom[39][103] = 16'hFFD2;
        rom[39][104] = 16'hFFFC;
        rom[39][105] = 16'h0002;
        rom[39][106] = 16'h000C;
        rom[39][107] = 16'hFFF9;
        rom[39][108] = 16'hFFD2;
        rom[39][109] = 16'hFFCD;
        rom[39][110] = 16'h0023;
        rom[39][111] = 16'h0004;
        rom[39][112] = 16'h0015;
        rom[39][113] = 16'h0005;
        rom[39][114] = 16'hFFCD;
        rom[39][115] = 16'hFFEF;
        rom[39][116] = 16'h0007;
        rom[39][117] = 16'h0030;
        rom[39][118] = 16'h000B;
        rom[39][119] = 16'hFFE4;
        rom[39][120] = 16'hFFF4;
        rom[39][121] = 16'hFFD2;
        rom[39][122] = 16'h001D;
        rom[39][123] = 16'h001D;
        rom[39][124] = 16'h0015;
        rom[39][125] = 16'h0004;
        rom[39][126] = 16'h0016;
        rom[39][127] = 16'h0024;
        rom[40][0] = 16'hFFD7;
        rom[40][1] = 16'h000F;
        rom[40][2] = 16'h0009;
        rom[40][3] = 16'hFFED;
        rom[40][4] = 16'hFFE1;
        rom[40][5] = 16'h0008;
        rom[40][6] = 16'hFFFC;
        rom[40][7] = 16'h001C;
        rom[40][8] = 16'hFFE6;
        rom[40][9] = 16'h0017;
        rom[40][10] = 16'hFFE1;
        rom[40][11] = 16'h0000;
        rom[40][12] = 16'h0013;
        rom[40][13] = 16'h0002;
        rom[40][14] = 16'h0001;
        rom[40][15] = 16'h0033;
        rom[40][16] = 16'hFFEB;
        rom[40][17] = 16'hFFD5;
        rom[40][18] = 16'h0015;
        rom[40][19] = 16'hFFE3;
        rom[40][20] = 16'h0018;
        rom[40][21] = 16'h000B;
        rom[40][22] = 16'hFFEF;
        rom[40][23] = 16'hFFDF;
        rom[40][24] = 16'h0011;
        rom[40][25] = 16'h0016;
        rom[40][26] = 16'h0007;
        rom[40][27] = 16'hFFEA;
        rom[40][28] = 16'hFFCB;
        rom[40][29] = 16'h0007;
        rom[40][30] = 16'hFFF4;
        rom[40][31] = 16'h0007;
        rom[40][32] = 16'h0004;
        rom[40][33] = 16'h0018;
        rom[40][34] = 16'hFFBB;
        rom[40][35] = 16'h0018;
        rom[40][36] = 16'h0012;
        rom[40][37] = 16'hFFCA;
        rom[40][38] = 16'hFFF6;
        rom[40][39] = 16'hFFCD;
        rom[40][40] = 16'h0009;
        rom[40][41] = 16'hFFF4;
        rom[40][42] = 16'h001B;
        rom[40][43] = 16'hFFC6;
        rom[40][44] = 16'h0019;
        rom[40][45] = 16'h000F;
        rom[40][46] = 16'hFFEC;
        rom[40][47] = 16'h0004;
        rom[40][48] = 16'h0015;
        rom[40][49] = 16'h0041;
        rom[40][50] = 16'hFFE1;
        rom[40][51] = 16'hFFEC;
        rom[40][52] = 16'hFFEF;
        rom[40][53] = 16'h001D;
        rom[40][54] = 16'hFFEF;
        rom[40][55] = 16'h0032;
        rom[40][56] = 16'h0030;
        rom[40][57] = 16'hFFDA;
        rom[40][58] = 16'hFFDA;
        rom[40][59] = 16'h000C;
        rom[40][60] = 16'hFFE7;
        rom[40][61] = 16'h0018;
        rom[40][62] = 16'h000C;
        rom[40][63] = 16'hFFE3;
        rom[40][64] = 16'hFFD5;
        rom[40][65] = 16'hFFEB;
        rom[40][66] = 16'hFFFE;
        rom[40][67] = 16'h000C;
        rom[40][68] = 16'hFFFC;
        rom[40][69] = 16'h002A;
        rom[40][70] = 16'h0020;
        rom[40][71] = 16'h0000;
        rom[40][72] = 16'h0010;
        rom[40][73] = 16'h003E;
        rom[40][74] = 16'hFFFE;
        rom[40][75] = 16'h0001;
        rom[40][76] = 16'h0000;
        rom[40][77] = 16'hFFE5;
        rom[40][78] = 16'hFFCF;
        rom[40][79] = 16'h000E;
        rom[40][80] = 16'hFFFB;
        rom[40][81] = 16'hFFE5;
        rom[40][82] = 16'hFFFE;
        rom[40][83] = 16'h004A;
        rom[40][84] = 16'h000C;
        rom[40][85] = 16'hFFF8;
        rom[40][86] = 16'h001F;
        rom[40][87] = 16'hFFD7;
        rom[40][88] = 16'hFFE5;
        rom[40][89] = 16'hFFF2;
        rom[40][90] = 16'hFFF6;
        rom[40][91] = 16'hFFE3;
        rom[40][92] = 16'hFFE4;
        rom[40][93] = 16'hFFD7;
        rom[40][94] = 16'hFFF2;
        rom[40][95] = 16'hFFA3;
        rom[40][96] = 16'hFFEF;
        rom[40][97] = 16'hFFDD;
        rom[40][98] = 16'hFFB4;
        rom[40][99] = 16'hFFC9;
        rom[40][100] = 16'hFFE8;
        rom[40][101] = 16'hFFED;
        rom[40][102] = 16'hFFBD;
        rom[40][103] = 16'hFFA3;
        rom[40][104] = 16'hFFF9;
        rom[40][105] = 16'hFFF1;
        rom[40][106] = 16'hFFE1;
        rom[40][107] = 16'h0025;
        rom[40][108] = 16'hFFF4;
        rom[40][109] = 16'h0002;
        rom[40][110] = 16'h0006;
        rom[40][111] = 16'h0006;
        rom[40][112] = 16'hFFD7;
        rom[40][113] = 16'hFFC8;
        rom[40][114] = 16'hFFC1;
        rom[40][115] = 16'hFFF0;
        rom[40][116] = 16'hFFC7;
        rom[40][117] = 16'h000B;
        rom[40][118] = 16'hFFE6;
        rom[40][119] = 16'hFFF9;
        rom[40][120] = 16'h0029;
        rom[40][121] = 16'hFFEE;
        rom[40][122] = 16'h000C;
        rom[40][123] = 16'hFFCE;
        rom[40][124] = 16'hFFEA;
        rom[40][125] = 16'hFFE2;
        rom[40][126] = 16'hFFCB;
        rom[40][127] = 16'h0004;
        rom[41][0] = 16'h0014;
        rom[41][1] = 16'hFFEF;
        rom[41][2] = 16'hFFA1;
        rom[41][3] = 16'h002C;
        rom[41][4] = 16'h002E;
        rom[41][5] = 16'hFFF7;
        rom[41][6] = 16'hFFD0;
        rom[41][7] = 16'hFFD9;
        rom[41][8] = 16'h0013;
        rom[41][9] = 16'hFFF8;
        rom[41][10] = 16'hFFEA;
        rom[41][11] = 16'hFFAB;
        rom[41][12] = 16'h0014;
        rom[41][13] = 16'hFFFB;
        rom[41][14] = 16'hFFF0;
        rom[41][15] = 16'hFFF8;
        rom[41][16] = 16'hFFCE;
        rom[41][17] = 16'hFFD7;
        rom[41][18] = 16'hFFC1;
        rom[41][19] = 16'hFFC3;
        rom[41][20] = 16'h0019;
        rom[41][21] = 16'hFFCF;
        rom[41][22] = 16'h0000;
        rom[41][23] = 16'hFFCB;
        rom[41][24] = 16'hFFD7;
        rom[41][25] = 16'h0003;
        rom[41][26] = 16'hFFA6;
        rom[41][27] = 16'h0017;
        rom[41][28] = 16'h0002;
        rom[41][29] = 16'h0007;
        rom[41][30] = 16'hFFD5;
        rom[41][31] = 16'h0012;
        rom[41][32] = 16'hFFF9;
        rom[41][33] = 16'hFFC2;
        rom[41][34] = 16'h0032;
        rom[41][35] = 16'h0032;
        rom[41][36] = 16'hFFEE;
        rom[41][37] = 16'h0011;
        rom[41][38] = 16'hFFEF;
        rom[41][39] = 16'h001E;
        rom[41][40] = 16'h000C;
        rom[41][41] = 16'hFFFD;
        rom[41][42] = 16'hFFFD;
        rom[41][43] = 16'h0012;
        rom[41][44] = 16'hFFF7;
        rom[41][45] = 16'hFFFC;
        rom[41][46] = 16'hFFD4;
        rom[41][47] = 16'h001C;
        rom[41][48] = 16'h0016;
        rom[41][49] = 16'hFFFB;
        rom[41][50] = 16'hFFED;
        rom[41][51] = 16'h001A;
        rom[41][52] = 16'hFFEE;
        rom[41][53] = 16'hFFEB;
        rom[41][54] = 16'hFFE1;
        rom[41][55] = 16'hFFEB;
        rom[41][56] = 16'hFFFD;
        rom[41][57] = 16'h002C;
        rom[41][58] = 16'hFFFC;
        rom[41][59] = 16'hFFCD;
        rom[41][60] = 16'hFFE0;
        rom[41][61] = 16'h0011;
        rom[41][62] = 16'hFFFF;
        rom[41][63] = 16'h0028;
        rom[41][64] = 16'h001F;
        rom[41][65] = 16'hFFBA;
        rom[41][66] = 16'hFFFB;
        rom[41][67] = 16'hFFFE;
        rom[41][68] = 16'hFFF8;
        rom[41][69] = 16'hFFFF;
        rom[41][70] = 16'hFFD6;
        rom[41][71] = 16'hFFD9;
        rom[41][72] = 16'hFFF9;
        rom[41][73] = 16'hFFF8;
        rom[41][74] = 16'h0010;
        rom[41][75] = 16'hFFBA;
        rom[41][76] = 16'hFFE2;
        rom[41][77] = 16'hFFDF;
        rom[41][78] = 16'hFFDD;
        rom[41][79] = 16'h001F;
        rom[41][80] = 16'hFFEB;
        rom[41][81] = 16'h001A;
        rom[41][82] = 16'hFFF6;
        rom[41][83] = 16'hFFED;
        rom[41][84] = 16'hFFE2;
        rom[41][85] = 16'h0009;
        rom[41][86] = 16'h0004;
        rom[41][87] = 16'hFFF4;
        rom[41][88] = 16'hFFD3;
        rom[41][89] = 16'h0024;
        rom[41][90] = 16'h0016;
        rom[41][91] = 16'h0007;
        rom[41][92] = 16'hFFE8;
        rom[41][93] = 16'h001B;
        rom[41][94] = 16'hFFC8;
        rom[41][95] = 16'h001A;
        rom[41][96] = 16'h0010;
        rom[41][97] = 16'h0006;
        rom[41][98] = 16'h0002;
        rom[41][99] = 16'h000B;
        rom[41][100] = 16'hFFF4;
        rom[41][101] = 16'h0011;
        rom[41][102] = 16'h0004;
        rom[41][103] = 16'h0011;
        rom[41][104] = 16'h0001;
        rom[41][105] = 16'h0016;
        rom[41][106] = 16'h0014;
        rom[41][107] = 16'hFFFB;
        rom[41][108] = 16'hFFAD;
        rom[41][109] = 16'h002D;
        rom[41][110] = 16'h0007;
        rom[41][111] = 16'hFFF9;
        rom[41][112] = 16'hFFE5;
        rom[41][113] = 16'hFFEA;
        rom[41][114] = 16'h000E;
        rom[41][115] = 16'hFFD5;
        rom[41][116] = 16'hFFCF;
        rom[41][117] = 16'hFFD5;
        rom[41][118] = 16'hFFF4;
        rom[41][119] = 16'hFFEC;
        rom[41][120] = 16'hFFE0;
        rom[41][121] = 16'hFFFD;
        rom[41][122] = 16'hFFAA;
        rom[41][123] = 16'h0014;
        rom[41][124] = 16'hFFDD;
        rom[41][125] = 16'h0014;
        rom[41][126] = 16'h0020;
        rom[41][127] = 16'h0005;
        rom[42][0] = 16'h0006;
        rom[42][1] = 16'hFFF2;
        rom[42][2] = 16'hFFE9;
        rom[42][3] = 16'hFFEC;
        rom[42][4] = 16'h0019;
        rom[42][5] = 16'hFFFB;
        rom[42][6] = 16'hFFC8;
        rom[42][7] = 16'h0024;
        rom[42][8] = 16'h0038;
        rom[42][9] = 16'h001E;
        rom[42][10] = 16'h0015;
        rom[42][11] = 16'h0027;
        rom[42][12] = 16'h0006;
        rom[42][13] = 16'h002A;
        rom[42][14] = 16'h0007;
        rom[42][15] = 16'h0007;
        rom[42][16] = 16'h001F;
        rom[42][17] = 16'hFFF9;
        rom[42][18] = 16'h0033;
        rom[42][19] = 16'h000E;
        rom[42][20] = 16'hFFFE;
        rom[42][21] = 16'h0004;
        rom[42][22] = 16'h002A;
        rom[42][23] = 16'hFFD7;
        rom[42][24] = 16'hFFDC;
        rom[42][25] = 16'hFFFE;
        rom[42][26] = 16'h0031;
        rom[42][27] = 16'hFFEE;
        rom[42][28] = 16'hFFE5;
        rom[42][29] = 16'hFFF8;
        rom[42][30] = 16'h0022;
        rom[42][31] = 16'h0037;
        rom[42][32] = 16'h002F;
        rom[42][33] = 16'h0011;
        rom[42][34] = 16'h0046;
        rom[42][35] = 16'h0004;
        rom[42][36] = 16'h0018;
        rom[42][37] = 16'hFFF9;
        rom[42][38] = 16'h0004;
        rom[42][39] = 16'hFFB5;
        rom[42][40] = 16'hFFF4;
        rom[42][41] = 16'hFFE8;
        rom[42][42] = 16'h0018;
        rom[42][43] = 16'hFFDC;
        rom[42][44] = 16'h0021;
        rom[42][45] = 16'h000B;
        rom[42][46] = 16'h0007;
        rom[42][47] = 16'hFFD2;
        rom[42][48] = 16'h001B;
        rom[42][49] = 16'hFFFB;
        rom[42][50] = 16'hFFC0;
        rom[42][51] = 16'hFFE8;
        rom[42][52] = 16'hFFF8;
        rom[42][53] = 16'hFFE7;
        rom[42][54] = 16'hFFF4;
        rom[42][55] = 16'hFFD9;
        rom[42][56] = 16'h0011;
        rom[42][57] = 16'hFFE0;
        rom[42][58] = 16'hFFE8;
        rom[42][59] = 16'h0041;
        rom[42][60] = 16'h0034;
        rom[42][61] = 16'h0011;
        rom[42][62] = 16'hFFB5;
        rom[42][63] = 16'hFFE7;
        rom[42][64] = 16'hFFE5;
        rom[42][65] = 16'h001F;
        rom[42][66] = 16'hFFE9;
        rom[42][67] = 16'h0027;
        rom[42][68] = 16'hFFC1;
        rom[42][69] = 16'h000C;
        rom[42][70] = 16'h0014;
        rom[42][71] = 16'h000B;
        rom[42][72] = 16'h002C;
        rom[42][73] = 16'h0004;
        rom[42][74] = 16'hFFEF;
        rom[42][75] = 16'hFFE2;
        rom[42][76] = 16'hFFFE;
        rom[42][77] = 16'h001B;
        rom[42][78] = 16'hFFE3;
        rom[42][79] = 16'h0025;
        rom[42][80] = 16'hFFFA;
        rom[42][81] = 16'hFFCC;
        rom[42][82] = 16'h001E;
        rom[42][83] = 16'h0015;
        rom[42][84] = 16'h0024;
        rom[42][85] = 16'hFFFB;
        rom[42][86] = 16'hFFFC;
        rom[42][87] = 16'h0019;
        rom[42][88] = 16'hFFD7;
        rom[42][89] = 16'hFFB4;
        rom[42][90] = 16'hFFFB;
        rom[42][91] = 16'h000E;
        rom[42][92] = 16'hFFE8;
        rom[42][93] = 16'h002C;
        rom[42][94] = 16'hFFDC;
        rom[42][95] = 16'hFFF1;
        rom[42][96] = 16'hFFEC;
        rom[42][97] = 16'hFFF7;
        rom[42][98] = 16'hFFDA;
        rom[42][99] = 16'h0012;
        rom[42][100] = 16'hFFC1;
        rom[42][101] = 16'h0012;
        rom[42][102] = 16'hFFEA;
        rom[42][103] = 16'hFFDC;
        rom[42][104] = 16'hFFEB;
        rom[42][105] = 16'h0009;
        rom[42][106] = 16'hFFFE;
        rom[42][107] = 16'h0010;
        rom[42][108] = 16'h0025;
        rom[42][109] = 16'hFFE4;
        rom[42][110] = 16'h0023;
        rom[42][111] = 16'hFFEA;
        rom[42][112] = 16'hFFCC;
        rom[42][113] = 16'hFFC2;
        rom[42][114] = 16'hFFDC;
        rom[42][115] = 16'hFFF7;
        rom[42][116] = 16'h0014;
        rom[42][117] = 16'hFFF2;
        rom[42][118] = 16'hFFD7;
        rom[42][119] = 16'hFFF3;
        rom[42][120] = 16'h0032;
        rom[42][121] = 16'hFFD2;
        rom[42][122] = 16'h0007;
        rom[42][123] = 16'h0018;
        rom[42][124] = 16'h0003;
        rom[42][125] = 16'hFFF8;
        rom[42][126] = 16'h0008;
        rom[42][127] = 16'h0024;
        rom[43][0] = 16'h0024;
        rom[43][1] = 16'hFFF3;
        rom[43][2] = 16'hFFE8;
        rom[43][3] = 16'h000D;
        rom[43][4] = 16'hFFF1;
        rom[43][5] = 16'hFFB0;
        rom[43][6] = 16'hFFB3;
        rom[43][7] = 16'h000E;
        rom[43][8] = 16'h0006;
        rom[43][9] = 16'hFFF2;
        rom[43][10] = 16'hFFD0;
        rom[43][11] = 16'hFFEA;
        rom[43][12] = 16'hFFEE;
        rom[43][13] = 16'h0023;
        rom[43][14] = 16'h001B;
        rom[43][15] = 16'h0012;
        rom[43][16] = 16'h0017;
        rom[43][17] = 16'hFFEE;
        rom[43][18] = 16'hFFE5;
        rom[43][19] = 16'hFFED;
        rom[43][20] = 16'hFFEB;
        rom[43][21] = 16'hFFFB;
        rom[43][22] = 16'hFFEA;
        rom[43][23] = 16'hFFEE;
        rom[43][24] = 16'h0039;
        rom[43][25] = 16'hFFDB;
        rom[43][26] = 16'h0001;
        rom[43][27] = 16'hFFFB;
        rom[43][28] = 16'h0002;
        rom[43][29] = 16'hFFF7;
        rom[43][30] = 16'h0013;
        rom[43][31] = 16'h0037;
        rom[43][32] = 16'hFFC9;
        rom[43][33] = 16'h0019;
        rom[43][34] = 16'h0023;
        rom[43][35] = 16'hFFFC;
        rom[43][36] = 16'hFFE7;
        rom[43][37] = 16'h0010;
        rom[43][38] = 16'h0027;
        rom[43][39] = 16'h001F;
        rom[43][40] = 16'hFFC2;
        rom[43][41] = 16'hFFED;
        rom[43][42] = 16'h0008;
        rom[43][43] = 16'hFFF4;
        rom[43][44] = 16'h001E;
        rom[43][45] = 16'h000A;
        rom[43][46] = 16'hFFE3;
        rom[43][47] = 16'hFFB0;
        rom[43][48] = 16'hFFF8;
        rom[43][49] = 16'hFFC2;
        rom[43][50] = 16'h000B;
        rom[43][51] = 16'hFFBB;
        rom[43][52] = 16'h0016;
        rom[43][53] = 16'hFFD9;
        rom[43][54] = 16'h002A;
        rom[43][55] = 16'hFFED;
        rom[43][56] = 16'h0002;
        rom[43][57] = 16'hFFE1;
        rom[43][58] = 16'h000D;
        rom[43][59] = 16'hFFFA;
        rom[43][60] = 16'hFFF9;
        rom[43][61] = 16'hFFDA;
        rom[43][62] = 16'hFFFC;
        rom[43][63] = 16'hFFBA;
        rom[43][64] = 16'hFFEF;
        rom[43][65] = 16'h0029;
        rom[43][66] = 16'hFFCD;
        rom[43][67] = 16'hFFC4;
        rom[43][68] = 16'h0002;
        rom[43][69] = 16'hFFAF;
        rom[43][70] = 16'h0009;
        rom[43][71] = 16'hFFFE;
        rom[43][72] = 16'h0016;
        rom[43][73] = 16'hFFDE;
        rom[43][74] = 16'hFFF4;
        rom[43][75] = 16'h0038;
        rom[43][76] = 16'h0027;
        rom[43][77] = 16'hFFF5;
        rom[43][78] = 16'h0008;
        rom[43][79] = 16'h001D;
        rom[43][80] = 16'hFFD0;
        rom[43][81] = 16'hFFED;
        rom[43][82] = 16'hFFBB;
        rom[43][83] = 16'h0004;
        rom[43][84] = 16'h000C;
        rom[43][85] = 16'h0011;
        rom[43][86] = 16'h0002;
        rom[43][87] = 16'h0027;
        rom[43][88] = 16'hFFCB;
        rom[43][89] = 16'h001D;
        rom[43][90] = 16'hFFC8;
        rom[43][91] = 16'hFFFB;
        rom[43][92] = 16'hFFFE;
        rom[43][93] = 16'hFFF7;
        rom[43][94] = 16'hFFFD;
        rom[43][95] = 16'h001B;
        rom[43][96] = 16'h000E;
        rom[43][97] = 16'hFFDD;
        rom[43][98] = 16'hFFD3;
        rom[43][99] = 16'h0018;
        rom[43][100] = 16'h000B;
        rom[43][101] = 16'hFFD7;
        rom[43][102] = 16'hFFCD;
        rom[43][103] = 16'h000E;
        rom[43][104] = 16'hFFD6;
        rom[43][105] = 16'h0038;
        rom[43][106] = 16'hFFD9;
        rom[43][107] = 16'h001C;
        rom[43][108] = 16'hFFF0;
        rom[43][109] = 16'hFFF9;
        rom[43][110] = 16'hFFCA;
        rom[43][111] = 16'hFFDE;
        rom[43][112] = 16'hFFE0;
        rom[43][113] = 16'hFFEA;
        rom[43][114] = 16'hFFE1;
        rom[43][115] = 16'h001F;
        rom[43][116] = 16'h0024;
        rom[43][117] = 16'hFFFD;
        rom[43][118] = 16'hFFA2;
        rom[43][119] = 16'h0007;
        rom[43][120] = 16'h001F;
        rom[43][121] = 16'h0006;
        rom[43][122] = 16'h0017;
        rom[43][123] = 16'h000B;
        rom[43][124] = 16'h001F;
        rom[43][125] = 16'hFFD4;
        rom[43][126] = 16'h0020;
        rom[43][127] = 16'hFFF4;
        rom[44][0] = 16'hFFF4;
        rom[44][1] = 16'hFFE1;
        rom[44][2] = 16'h0011;
        rom[44][3] = 16'h000C;
        rom[44][4] = 16'hFFF5;
        rom[44][5] = 16'h0022;
        rom[44][6] = 16'hFFD2;
        rom[44][7] = 16'hFFC2;
        rom[44][8] = 16'h0024;
        rom[44][9] = 16'h002F;
        rom[44][10] = 16'hFFEF;
        rom[44][11] = 16'h0008;
        rom[44][12] = 16'hFFFC;
        rom[44][13] = 16'hFFF6;
        rom[44][14] = 16'hFFFE;
        rom[44][15] = 16'h0013;
        rom[44][16] = 16'hFFF0;
        rom[44][17] = 16'hFFF9;
        rom[44][18] = 16'hFFC3;
        rom[44][19] = 16'hFFE5;
        rom[44][20] = 16'hFFDF;
        rom[44][21] = 16'h0007;
        rom[44][22] = 16'hFFDD;
        rom[44][23] = 16'hFFBA;
        rom[44][24] = 16'h0012;
        rom[44][25] = 16'h0009;
        rom[44][26] = 16'hFFE7;
        rom[44][27] = 16'h0020;
        rom[44][28] = 16'hFFFF;
        rom[44][29] = 16'hFFD9;
        rom[44][30] = 16'hFFF7;
        rom[44][31] = 16'hFFF3;
        rom[44][32] = 16'hFFFE;
        rom[44][33] = 16'hFFCA;
        rom[44][34] = 16'hFFF6;
        rom[44][35] = 16'h0002;
        rom[44][36] = 16'hFFBB;
        rom[44][37] = 16'hFFEE;
        rom[44][38] = 16'hFFE4;
        rom[44][39] = 16'hFFF3;
        rom[44][40] = 16'h0027;
        rom[44][41] = 16'hFFF4;
        rom[44][42] = 16'hFFC4;
        rom[44][43] = 16'hFFE0;
        rom[44][44] = 16'hFFE0;
        rom[44][45] = 16'h000F;
        rom[44][46] = 16'hFFE1;
        rom[44][47] = 16'hFFEA;
        rom[44][48] = 16'hFFE6;
        rom[44][49] = 16'hFFE9;
        rom[44][50] = 16'h0009;
        rom[44][51] = 16'h000B;
        rom[44][52] = 16'h0011;
        rom[44][53] = 16'h0032;
        rom[44][54] = 16'h0007;
        rom[44][55] = 16'h0029;
        rom[44][56] = 16'h0019;
        rom[44][57] = 16'h0012;
        rom[44][58] = 16'hFFCF;
        rom[44][59] = 16'hFFF5;
        rom[44][60] = 16'hFFE5;
        rom[44][61] = 16'hFFDB;
        rom[44][62] = 16'h0024;
        rom[44][63] = 16'hFFDD;
        rom[44][64] = 16'hFFE5;
        rom[44][65] = 16'hFFBA;
        rom[44][66] = 16'h000C;
        rom[44][67] = 16'h0016;
        rom[44][68] = 16'h0018;
        rom[44][69] = 16'hFFFB;
        rom[44][70] = 16'h0014;
        rom[44][71] = 16'hFFF4;
        rom[44][72] = 16'h0017;
        rom[44][73] = 16'h0017;
        rom[44][74] = 16'hFFE3;
        rom[44][75] = 16'h000B;
        rom[44][76] = 16'h001E;
        rom[44][77] = 16'h0001;
        rom[44][78] = 16'hFFF2;
        rom[44][79] = 16'h0006;
        rom[44][80] = 16'h0007;
        rom[44][81] = 16'hFFF9;
        rom[44][82] = 16'hFFFA;
        rom[44][83] = 16'hFFE5;
        rom[44][84] = 16'hFFB2;
        rom[44][85] = 16'h000E;
        rom[44][86] = 16'h0019;
        rom[44][87] = 16'hFFF4;
        rom[44][88] = 16'hFFD2;
        rom[44][89] = 16'h0002;
        rom[44][90] = 16'hFFF9;
        rom[44][91] = 16'hFFE6;
        rom[44][92] = 16'hFFF5;
        rom[44][93] = 16'hFFEE;
        rom[44][94] = 16'hFFF9;
        rom[44][95] = 16'hFFB8;
        rom[44][96] = 16'hFFED;
        rom[44][97] = 16'hFFF4;
        rom[44][98] = 16'hFFFE;
        rom[44][99] = 16'hFFCD;
        rom[44][100] = 16'hFFF3;
        rom[44][101] = 16'hFFF9;
        rom[44][102] = 16'h000C;
        rom[44][103] = 16'hFFF8;
        rom[44][104] = 16'h0016;
        rom[44][105] = 16'hFFEA;
        rom[44][106] = 16'h0004;
        rom[44][107] = 16'h0016;
        rom[44][108] = 16'h0012;
        rom[44][109] = 16'h0021;
        rom[44][110] = 16'hFFDB;
        rom[44][111] = 16'h0002;
        rom[44][112] = 16'hFFFE;
        rom[44][113] = 16'hFFFA;
        rom[44][114] = 16'h0001;
        rom[44][115] = 16'h0007;
        rom[44][116] = 16'hFFC8;
        rom[44][117] = 16'h0001;
        rom[44][118] = 16'hFFED;
        rom[44][119] = 16'hFFEF;
        rom[44][120] = 16'hFFEC;
        rom[44][121] = 16'h0020;
        rom[44][122] = 16'h0004;
        rom[44][123] = 16'h0002;
        rom[44][124] = 16'hFFDD;
        rom[44][125] = 16'h0024;
        rom[44][126] = 16'h001F;
        rom[44][127] = 16'hFFF5;
        rom[45][0] = 16'h0009;
        rom[45][1] = 16'h002E;
        rom[45][2] = 16'hFFF5;
        rom[45][3] = 16'h001F;
        rom[45][4] = 16'h0025;
        rom[45][5] = 16'h0031;
        rom[45][6] = 16'h0006;
        rom[45][7] = 16'h0022;
        rom[45][8] = 16'hFFFF;
        rom[45][9] = 16'hFFC3;
        rom[45][10] = 16'hFFB7;
        rom[45][11] = 16'h0002;
        rom[45][12] = 16'hFFC3;
        rom[45][13] = 16'hFFAA;
        rom[45][14] = 16'hFFF9;
        rom[45][15] = 16'h0015;
        rom[45][16] = 16'h0023;
        rom[45][17] = 16'hFFF9;
        rom[45][18] = 16'hFFD3;
        rom[45][19] = 16'hFFE0;
        rom[45][20] = 16'hFFF3;
        rom[45][21] = 16'hFFFA;
        rom[45][22] = 16'hFFC7;
        rom[45][23] = 16'hFFDD;
        rom[45][24] = 16'hFFFF;
        rom[45][25] = 16'hFFD6;
        rom[45][26] = 16'h0013;
        rom[45][27] = 16'hFFE9;
        rom[45][28] = 16'h000C;
        rom[45][29] = 16'hFFCF;
        rom[45][30] = 16'h0007;
        rom[45][31] = 16'h0006;
        rom[45][32] = 16'h0004;
        rom[45][33] = 16'h0019;
        rom[45][34] = 16'hFFD2;
        rom[45][35] = 16'h0011;
        rom[45][36] = 16'hFFEC;
        rom[45][37] = 16'h000D;
        rom[45][38] = 16'hFFF7;
        rom[45][39] = 16'hFFE7;
        rom[45][40] = 16'hFFC2;
        rom[45][41] = 16'hFFBF;
        rom[45][42] = 16'hFF97;
        rom[45][43] = 16'h0012;
        rom[45][44] = 16'hFFDB;
        rom[45][45] = 16'h0003;
        rom[45][46] = 16'h0010;
        rom[45][47] = 16'hFFF3;
        rom[45][48] = 16'hFFF9;
        rom[45][49] = 16'h0005;
        rom[45][50] = 16'h001A;
        rom[45][51] = 16'h0001;
        rom[45][52] = 16'h0016;
        rom[45][53] = 16'h0000;
        rom[45][54] = 16'h0028;
        rom[45][55] = 16'hFFDE;
        rom[45][56] = 16'hFFDC;
        rom[45][57] = 16'h001F;
        rom[45][58] = 16'h0002;
        rom[45][59] = 16'hFFEE;
        rom[45][60] = 16'h000E;
        rom[45][61] = 16'hFFE5;
        rom[45][62] = 16'h0017;
        rom[45][63] = 16'h001E;
        rom[45][64] = 16'hFFF8;
        rom[45][65] = 16'h0018;
        rom[45][66] = 16'h001F;
        rom[45][67] = 16'h0022;
        rom[45][68] = 16'hFFE4;
        rom[45][69] = 16'h0008;
        rom[45][70] = 16'h001B;
        rom[45][71] = 16'h002C;
        rom[45][72] = 16'hFFC2;
        rom[45][73] = 16'hFFFA;
        rom[45][74] = 16'hFFFA;
        rom[45][75] = 16'h000E;
        rom[45][76] = 16'hFFEB;
        rom[45][77] = 16'hFFF8;
        rom[45][78] = 16'h000D;
        rom[45][79] = 16'hFFEA;
        rom[45][80] = 16'h0025;
        rom[45][81] = 16'h0027;
        rom[45][82] = 16'h0032;
        rom[45][83] = 16'hFFD8;
        rom[45][84] = 16'hFFF2;
        rom[45][85] = 16'h001A;
        rom[45][86] = 16'hFFC9;
        rom[45][87] = 16'h000B;
        rom[45][88] = 16'hFFE5;
        rom[45][89] = 16'h0023;
        rom[45][90] = 16'h000B;
        rom[45][91] = 16'h0028;
        rom[45][92] = 16'h0025;
        rom[45][93] = 16'h0016;
        rom[45][94] = 16'h0011;
        rom[45][95] = 16'hFFFC;
        rom[45][96] = 16'hFFF6;
        rom[45][97] = 16'hFFF4;
        rom[45][98] = 16'hFFF7;
        rom[45][99] = 16'h0021;
        rom[45][100] = 16'hFFEC;
        rom[45][101] = 16'h0016;
        rom[45][102] = 16'h0023;
        rom[45][103] = 16'hFFFA;
        rom[45][104] = 16'hFFFC;
        rom[45][105] = 16'hFFE7;
        rom[45][106] = 16'hFFE1;
        rom[45][107] = 16'hFFE1;
        rom[45][108] = 16'hFFF7;
        rom[45][109] = 16'hFFFB;
        rom[45][110] = 16'h002B;
        rom[45][111] = 16'h0013;
        rom[45][112] = 16'h001F;
        rom[45][113] = 16'h0009;
        rom[45][114] = 16'h0011;
        rom[45][115] = 16'h0014;
        rom[45][116] = 16'h0033;
        rom[45][117] = 16'hFFDF;
        rom[45][118] = 16'h0014;
        rom[45][119] = 16'hFFFD;
        rom[45][120] = 16'hFFEE;
        rom[45][121] = 16'hFFE4;
        rom[45][122] = 16'hFFF9;
        rom[45][123] = 16'h001A;
        rom[45][124] = 16'h0038;
        rom[45][125] = 16'h0004;
        rom[45][126] = 16'h003D;
        rom[45][127] = 16'hFFDF;
        rom[46][0] = 16'hFFDD;
        rom[46][1] = 16'hFFEA;
        rom[46][2] = 16'h000B;
        rom[46][3] = 16'hFFDC;
        rom[46][4] = 16'h0001;
        rom[46][5] = 16'h0006;
        rom[46][6] = 16'hFFC4;
        rom[46][7] = 16'hFFC2;
        rom[46][8] = 16'hFFE5;
        rom[46][9] = 16'hFFF1;
        rom[46][10] = 16'hFFF1;
        rom[46][11] = 16'hFFE4;
        rom[46][12] = 16'hFFC3;
        rom[46][13] = 16'hFFD5;
        rom[46][14] = 16'h0050;
        rom[46][15] = 16'h0014;
        rom[46][16] = 16'hFFE1;
        rom[46][17] = 16'hFFF2;
        rom[46][18] = 16'hFFCC;
        rom[46][19] = 16'hFFDE;
        rom[46][20] = 16'hFFEA;
        rom[46][21] = 16'hFFF9;
        rom[46][22] = 16'hFFF7;
        rom[46][23] = 16'hFFDA;
        rom[46][24] = 16'h0017;
        rom[46][25] = 16'h0007;
        rom[46][26] = 16'h0011;
        rom[46][27] = 16'h0025;
        rom[46][28] = 16'h0020;
        rom[46][29] = 16'hFFFE;
        rom[46][30] = 16'h0010;
        rom[46][31] = 16'hFFFA;
        rom[46][32] = 16'hFFF9;
        rom[46][33] = 16'hFFE5;
        rom[46][34] = 16'hFFF4;
        rom[46][35] = 16'hFFFA;
        rom[46][36] = 16'hFFA6;
        rom[46][37] = 16'hFFCE;
        rom[46][38] = 16'hFFF9;
        rom[46][39] = 16'hFFDA;
        rom[46][40] = 16'hFFFB;
        rom[46][41] = 16'hFFDD;
        rom[46][42] = 16'hFFF3;
        rom[46][43] = 16'h0002;
        rom[46][44] = 16'h0001;
        rom[46][45] = 16'h0012;
        rom[46][46] = 16'hFFCD;
        rom[46][47] = 16'hFFD7;
        rom[46][48] = 16'hFFF2;
        rom[46][49] = 16'h0017;
        rom[46][50] = 16'h0006;
        rom[46][51] = 16'h001D;
        rom[46][52] = 16'h0028;
        rom[46][53] = 16'hFFF5;
        rom[46][54] = 16'h0006;
        rom[46][55] = 16'hFFF8;
        rom[46][56] = 16'h001E;
        rom[46][57] = 16'h001C;
        rom[46][58] = 16'hFFE5;
        rom[46][59] = 16'h001D;
        rom[46][60] = 16'hFFF8;
        rom[46][61] = 16'h0001;
        rom[46][62] = 16'hFFFD;
        rom[46][63] = 16'hFFF9;
        rom[46][64] = 16'hFFC8;
        rom[46][65] = 16'hFFE1;
        rom[46][66] = 16'h0014;
        rom[46][67] = 16'hFFEF;
        rom[46][68] = 16'h0010;
        rom[46][69] = 16'hFFF8;
        rom[46][70] = 16'h001A;
        rom[46][71] = 16'h0002;
        rom[46][72] = 16'hFFE4;
        rom[46][73] = 16'h000C;
        rom[46][74] = 16'hFFC3;
        rom[46][75] = 16'h001F;
        rom[46][76] = 16'h002D;
        rom[46][77] = 16'hFFFC;
        rom[46][78] = 16'hFFED;
        rom[46][79] = 16'h0005;
        rom[46][80] = 16'h0014;
        rom[46][81] = 16'hFFE5;
        rom[46][82] = 16'h0015;
        rom[46][83] = 16'hFFF6;
        rom[46][84] = 16'hFFDE;
        rom[46][85] = 16'hFFFF;
        rom[46][86] = 16'hFFF3;
        rom[46][87] = 16'h0000;
        rom[46][88] = 16'hFFF4;
        rom[46][89] = 16'h0025;
        rom[46][90] = 16'h0009;
        rom[46][91] = 16'h0019;
        rom[46][92] = 16'hFFED;
        rom[46][93] = 16'hFFEA;
        rom[46][94] = 16'hFFE1;
        rom[46][95] = 16'hFFCC;
        rom[46][96] = 16'h0020;
        rom[46][97] = 16'hFFEE;
        rom[46][98] = 16'hFFF5;
        rom[46][99] = 16'hFFCD;
        rom[46][100] = 16'hFFE8;
        rom[46][101] = 16'hFFF2;
        rom[46][102] = 16'hFFEE;
        rom[46][103] = 16'hFFF9;
        rom[46][104] = 16'h0007;
        rom[46][105] = 16'hFFD4;
        rom[46][106] = 16'h0014;
        rom[46][107] = 16'h0002;
        rom[46][108] = 16'h0010;
        rom[46][109] = 16'h0008;
        rom[46][110] = 16'h0012;
        rom[46][111] = 16'hFFF1;
        rom[46][112] = 16'h003E;
        rom[46][113] = 16'hFFDD;
        rom[46][114] = 16'h0019;
        rom[46][115] = 16'hFFEB;
        rom[46][116] = 16'hFFCA;
        rom[46][117] = 16'h0039;
        rom[46][118] = 16'h002A;
        rom[46][119] = 16'hFFE8;
        rom[46][120] = 16'hFFD7;
        rom[46][121] = 16'hFFF4;
        rom[46][122] = 16'h000E;
        rom[46][123] = 16'h0001;
        rom[46][124] = 16'h0024;
        rom[46][125] = 16'h0024;
        rom[46][126] = 16'h0019;
        rom[46][127] = 16'hFFFF;
        rom[47][0] = 16'h0051;
        rom[47][1] = 16'hFFF7;
        rom[47][2] = 16'h0010;
        rom[47][3] = 16'h0018;
        rom[47][4] = 16'h0005;
        rom[47][5] = 16'hFFEF;
        rom[47][6] = 16'hFFD2;
        rom[47][7] = 16'hFFF3;
        rom[47][8] = 16'h0004;
        rom[47][9] = 16'h0016;
        rom[47][10] = 16'hFFD6;
        rom[47][11] = 16'hFFEA;
        rom[47][12] = 16'hFFEF;
        rom[47][13] = 16'hFFD7;
        rom[47][14] = 16'hFFE5;
        rom[47][15] = 16'h0002;
        rom[47][16] = 16'hFFDD;
        rom[47][17] = 16'hFFF0;
        rom[47][18] = 16'h0019;
        rom[47][19] = 16'hFFF3;
        rom[47][20] = 16'hFFFA;
        rom[47][21] = 16'h004F;
        rom[47][22] = 16'hFFBC;
        rom[47][23] = 16'h0009;
        rom[47][24] = 16'h0024;
        rom[47][25] = 16'hFFDD;
        rom[47][26] = 16'h001B;
        rom[47][27] = 16'hFFFD;
        rom[47][28] = 16'hFFED;
        rom[47][29] = 16'hFFDD;
        rom[47][30] = 16'hFFF8;
        rom[47][31] = 16'h002F;
        rom[47][32] = 16'hFFF5;
        rom[47][33] = 16'h0016;
        rom[47][34] = 16'hFFE9;
        rom[47][35] = 16'hFFC7;
        rom[47][36] = 16'hFFC3;
        rom[47][37] = 16'h0019;
        rom[47][38] = 16'hFFED;
        rom[47][39] = 16'hFFF7;
        rom[47][40] = 16'hFFCD;
        rom[47][41] = 16'h0056;
        rom[47][42] = 16'h0021;
        rom[47][43] = 16'h0012;
        rom[47][44] = 16'h000B;
        rom[47][45] = 16'hFFEE;
        rom[47][46] = 16'hFFDF;
        rom[47][47] = 16'hFFFE;
        rom[47][48] = 16'hFFFE;
        rom[47][49] = 16'hFFE8;
        rom[47][50] = 16'hFFD0;
        rom[47][51] = 16'h0008;
        rom[47][52] = 16'h0004;
        rom[47][53] = 16'h001B;
        rom[47][54] = 16'hFFFC;
        rom[47][55] = 16'hFFE0;
        rom[47][56] = 16'h0015;
        rom[47][57] = 16'h002B;
        rom[47][58] = 16'h0012;
        rom[47][59] = 16'hFFDA;
        rom[47][60] = 16'hFFB3;
        rom[47][61] = 16'h000C;
        rom[47][62] = 16'hFFA4;
        rom[47][63] = 16'h001B;
        rom[47][64] = 16'h0023;
        rom[47][65] = 16'h001F;
        rom[47][66] = 16'hFFF0;
        rom[47][67] = 16'h000B;
        rom[47][68] = 16'h0005;
        rom[47][69] = 16'hFFCA;
        rom[47][70] = 16'hFFEF;
        rom[47][71] = 16'h0003;
        rom[47][72] = 16'h0035;
        rom[47][73] = 16'hFFE5;
        rom[47][74] = 16'h002A;
        rom[47][75] = 16'h0024;
        rom[47][76] = 16'h0013;
        rom[47][77] = 16'hFFF5;
        rom[47][78] = 16'h001F;
        rom[47][79] = 16'h0024;
        rom[47][80] = 16'hFFC9;
        rom[47][81] = 16'hFFC6;
        rom[47][82] = 16'hFFF4;
        rom[47][83] = 16'hFFE2;
        rom[47][84] = 16'hFFDA;
        rom[47][85] = 16'h0008;
        rom[47][86] = 16'h001D;
        rom[47][87] = 16'hFFEE;
        rom[47][88] = 16'hFFF4;
        rom[47][89] = 16'h0009;
        rom[47][90] = 16'hFFF8;
        rom[47][91] = 16'h0016;
        rom[47][92] = 16'h000C;
        rom[47][93] = 16'hFFCC;
        rom[47][94] = 16'hFFF6;
        rom[47][95] = 16'hFFF9;
        rom[47][96] = 16'hFFE0;
        rom[47][97] = 16'hFFF7;
        rom[47][98] = 16'h0021;
        rom[47][99] = 16'hFFD2;
        rom[47][100] = 16'hFFF4;
        rom[47][101] = 16'h002B;
        rom[47][102] = 16'hFFC5;
        rom[47][103] = 16'hFFEA;
        rom[47][104] = 16'h0039;
        rom[47][105] = 16'h000E;
        rom[47][106] = 16'hFFFB;
        rom[47][107] = 16'hFFB6;
        rom[47][108] = 16'h0014;
        rom[47][109] = 16'hFFEF;
        rom[47][110] = 16'hFFE7;
        rom[47][111] = 16'hFFC3;
        rom[47][112] = 16'h0009;
        rom[47][113] = 16'h0000;
        rom[47][114] = 16'hFFCE;
        rom[47][115] = 16'hFFD1;
        rom[47][116] = 16'hFFD4;
        rom[47][117] = 16'hFFE1;
        rom[47][118] = 16'hFFED;
        rom[47][119] = 16'hFFE6;
        rom[47][120] = 16'h0021;
        rom[47][121] = 16'hFFDA;
        rom[47][122] = 16'hFFF9;
        rom[47][123] = 16'h0011;
        rom[47][124] = 16'hFFF0;
        rom[47][125] = 16'h0018;
        rom[47][126] = 16'hFFDA;
        rom[47][127] = 16'hFFEF;
        rom[48][0] = 16'h0014;
        rom[48][1] = 16'hFFFB;
        rom[48][2] = 16'hFFDF;
        rom[48][3] = 16'hFFEC;
        rom[48][4] = 16'h001F;
        rom[48][5] = 16'hFFED;
        rom[48][6] = 16'hFFBD;
        rom[48][7] = 16'hFFE6;
        rom[48][8] = 16'h0024;
        rom[48][9] = 16'h0004;
        rom[48][10] = 16'hFFBB;
        rom[48][11] = 16'h0011;
        rom[48][12] = 16'hFFE9;
        rom[48][13] = 16'hFFF4;
        rom[48][14] = 16'hFFDF;
        rom[48][15] = 16'hFFFE;
        rom[48][16] = 16'hFFEE;
        rom[48][17] = 16'hFFFE;
        rom[48][18] = 16'hFFFF;
        rom[48][19] = 16'h0007;
        rom[48][20] = 16'h0004;
        rom[48][21] = 16'h0007;
        rom[48][22] = 16'hFFDA;
        rom[48][23] = 16'h0002;
        rom[48][24] = 16'h0016;
        rom[48][25] = 16'hFFEA;
        rom[48][26] = 16'h0007;
        rom[48][27] = 16'hFFFF;
        rom[48][28] = 16'h0007;
        rom[48][29] = 16'h0023;
        rom[48][30] = 16'h0002;
        rom[48][31] = 16'hFFE5;
        rom[48][32] = 16'h001D;
        rom[48][33] = 16'h0003;
        rom[48][34] = 16'hFFD7;
        rom[48][35] = 16'h001B;
        rom[48][36] = 16'hFFE5;
        rom[48][37] = 16'h0024;
        rom[48][38] = 16'hFFD1;
        rom[48][39] = 16'h0006;
        rom[48][40] = 16'hFFE4;
        rom[48][41] = 16'hFFE5;
        rom[48][42] = 16'h000D;
        rom[48][43] = 16'h0037;
        rom[48][44] = 16'hFFFA;
        rom[48][45] = 16'h0006;
        rom[48][46] = 16'hFFF1;
        rom[48][47] = 16'h000D;
        rom[48][48] = 16'h0007;
        rom[48][49] = 16'h001D;
        rom[48][50] = 16'hFFB0;
        rom[48][51] = 16'hFFF2;
        rom[48][52] = 16'hFFB9;
        rom[48][53] = 16'h001C;
        rom[48][54] = 16'hFFC7;
        rom[48][55] = 16'h000F;
        rom[48][56] = 16'h0011;
        rom[48][57] = 16'hFFFB;
        rom[48][58] = 16'h0023;
        rom[48][59] = 16'hFFFB;
        rom[48][60] = 16'h0012;
        rom[48][61] = 16'h000D;
        rom[48][62] = 16'hFFD4;
        rom[48][63] = 16'hFFC6;
        rom[48][64] = 16'hFFCE;
        rom[48][65] = 16'hFFF3;
        rom[48][66] = 16'hFFDC;
        rom[48][67] = 16'hFFEF;
        rom[48][68] = 16'h0020;
        rom[48][69] = 16'h0001;
        rom[48][70] = 16'hFFDB;
        rom[48][71] = 16'hFFE0;
        rom[48][72] = 16'h0016;
        rom[48][73] = 16'hFFFD;
        rom[48][74] = 16'hFFEF;
        rom[48][75] = 16'hFFF3;
        rom[48][76] = 16'hFFE5;
        rom[48][77] = 16'hFFA3;
        rom[48][78] = 16'hFFE5;
        rom[48][79] = 16'h0002;
        rom[48][80] = 16'h0005;
        rom[48][81] = 16'hFFCB;
        rom[48][82] = 16'h000D;
        rom[48][83] = 16'hFFFD;
        rom[48][84] = 16'hFFC1;
        rom[48][85] = 16'hFFB9;
        rom[48][86] = 16'h0018;
        rom[48][87] = 16'hFFFC;
        rom[48][88] = 16'hFFD4;
        rom[48][89] = 16'hFFD7;
        rom[48][90] = 16'h0006;
        rom[48][91] = 16'h0006;
        rom[48][92] = 16'h0001;
        rom[48][93] = 16'h0020;
        rom[48][94] = 16'hFFE7;
        rom[48][95] = 16'hFFFB;
        rom[48][96] = 16'hFFEA;
        rom[48][97] = 16'h0011;
        rom[48][98] = 16'h0029;
        rom[48][99] = 16'h0009;
        rom[48][100] = 16'h0004;
        rom[48][101] = 16'hFFD5;
        rom[48][102] = 16'hFFFB;
        rom[48][103] = 16'h0011;
        rom[48][104] = 16'hFFCC;
        rom[48][105] = 16'hFFCC;
        rom[48][106] = 16'hFFD3;
        rom[48][107] = 16'h0001;
        rom[48][108] = 16'h0006;
        rom[48][109] = 16'h0000;
        rom[48][110] = 16'h0008;
        rom[48][111] = 16'hFFFC;
        rom[48][112] = 16'hFFFC;
        rom[48][113] = 16'hFFDA;
        rom[48][114] = 16'h0017;
        rom[48][115] = 16'hFFE6;
        rom[48][116] = 16'h0011;
        rom[48][117] = 16'hFFF4;
        rom[48][118] = 16'h0002;
        rom[48][119] = 16'hFFB9;
        rom[48][120] = 16'hFFFE;
        rom[48][121] = 16'h001B;
        rom[48][122] = 16'h0007;
        rom[48][123] = 16'h0008;
        rom[48][124] = 16'hFFC8;
        rom[48][125] = 16'hFFC1;
        rom[48][126] = 16'h0010;
        rom[48][127] = 16'h0011;
        rom[49][0] = 16'hFFE6;
        rom[49][1] = 16'hFFC2;
        rom[49][2] = 16'h001A;
        rom[49][3] = 16'hFFFF;
        rom[49][4] = 16'hFFF9;
        rom[49][5] = 16'hFFE6;
        rom[49][6] = 16'hFFED;
        rom[49][7] = 16'hFFEF;
        rom[49][8] = 16'hFFE1;
        rom[49][9] = 16'h0015;
        rom[49][10] = 16'hFFF3;
        rom[49][11] = 16'hFFFB;
        rom[49][12] = 16'h0008;
        rom[49][13] = 16'h0007;
        rom[49][14] = 16'h001F;
        rom[49][15] = 16'h0008;
        rom[49][16] = 16'h0008;
        rom[49][17] = 16'h001F;
        rom[49][18] = 16'h0011;
        rom[49][19] = 16'h0014;
        rom[49][20] = 16'hFFEC;
        rom[49][21] = 16'hFFD3;
        rom[49][22] = 16'h0000;
        rom[49][23] = 16'h0002;
        rom[49][24] = 16'h0017;
        rom[49][25] = 16'hFFE2;
        rom[49][26] = 16'h0016;
        rom[49][27] = 16'h000E;
        rom[49][28] = 16'h0016;
        rom[49][29] = 16'h000C;
        rom[49][30] = 16'h0011;
        rom[49][31] = 16'hFFC0;
        rom[49][32] = 16'h0002;
        rom[49][33] = 16'hFFFF;
        rom[49][34] = 16'hFFF6;
        rom[49][35] = 16'h0003;
        rom[49][36] = 16'hFFC5;
        rom[49][37] = 16'h0002;
        rom[49][38] = 16'hFFEF;
        rom[49][39] = 16'h0015;
        rom[49][40] = 16'h0012;
        rom[49][41] = 16'hFFEC;
        rom[49][42] = 16'hFFB8;
        rom[49][43] = 16'h0029;
        rom[49][44] = 16'h0007;
        rom[49][45] = 16'hFFE5;
        rom[49][46] = 16'hFFCF;
        rom[49][47] = 16'hFFEF;
        rom[49][48] = 16'hFFD7;
        rom[49][49] = 16'h0068;
        rom[49][50] = 16'hFFFB;
        rom[49][51] = 16'h0012;
        rom[49][52] = 16'hFFEF;
        rom[49][53] = 16'h0020;
        rom[49][54] = 16'hFFDD;
        rom[49][55] = 16'hFFBB;
        rom[49][56] = 16'hFFCD;
        rom[49][57] = 16'hFFC8;
        rom[49][58] = 16'hFFD3;
        rom[49][59] = 16'h0007;
        rom[49][60] = 16'h0030;
        rom[49][61] = 16'h0007;
        rom[49][62] = 16'hFFD7;
        rom[49][63] = 16'hFFE8;
        rom[49][64] = 16'h0007;
        rom[49][65] = 16'hFFF5;
        rom[49][66] = 16'hFFF6;
        rom[49][67] = 16'hFFEF;
        rom[49][68] = 16'hFFEF;
        rom[49][69] = 16'h0011;
        rom[49][70] = 16'hFFD4;
        rom[49][71] = 16'h0003;
        rom[49][72] = 16'hFFF6;
        rom[49][73] = 16'h000C;
        rom[49][74] = 16'hFFCC;
        rom[49][75] = 16'hFFFE;
        rom[49][76] = 16'h0004;
        rom[49][77] = 16'hFFF2;
        rom[49][78] = 16'hFFEF;
        rom[49][79] = 16'hFFD7;
        rom[49][80] = 16'hFFF3;
        rom[49][81] = 16'hFFC9;
        rom[49][82] = 16'hFFFC;
        rom[49][83] = 16'hFFFD;
        rom[49][84] = 16'h0023;
        rom[49][85] = 16'h000F;
        rom[49][86] = 16'h001B;
        rom[49][87] = 16'hFFE1;
        rom[49][88] = 16'h002B;
        rom[49][89] = 16'hFFE0;
        rom[49][90] = 16'h0010;
        rom[49][91] = 16'h0000;
        rom[49][92] = 16'h0007;
        rom[49][93] = 16'h0016;
        rom[49][94] = 16'hFFE5;
        rom[49][95] = 16'hFFD7;
        rom[49][96] = 16'hFFE8;
        rom[49][97] = 16'hFFBB;
        rom[49][98] = 16'h002B;
        rom[49][99] = 16'hFFB6;
        rom[49][100] = 16'hFFFE;
        rom[49][101] = 16'hFFDF;
        rom[49][102] = 16'hFFBB;
        rom[49][103] = 16'hFFDF;
        rom[49][104] = 16'hFFDC;
        rom[49][105] = 16'hFFF3;
        rom[49][106] = 16'hFFDB;
        rom[49][107] = 16'hFFE4;
        rom[49][108] = 16'hFFFC;
        rom[49][109] = 16'hFFD8;
        rom[49][110] = 16'h001F;
        rom[49][111] = 16'h001B;
        rom[49][112] = 16'h0005;
        rom[49][113] = 16'h000F;
        rom[49][114] = 16'h0023;
        rom[49][115] = 16'hFFC3;
        rom[49][116] = 16'hFFFE;
        rom[49][117] = 16'h0014;
        rom[49][118] = 16'hFFE1;
        rom[49][119] = 16'hFFF4;
        rom[49][120] = 16'h0010;
        rom[49][121] = 16'h0029;
        rom[49][122] = 16'hFFFF;
        rom[49][123] = 16'h0014;
        rom[49][124] = 16'hFFF8;
        rom[49][125] = 16'hFFEB;
        rom[49][126] = 16'h0020;
        rom[49][127] = 16'hFFF4;
        rom[50][0] = 16'hFFF8;
        rom[50][1] = 16'h0000;
        rom[50][2] = 16'hFFDC;
        rom[50][3] = 16'hFFEF;
        rom[50][4] = 16'h0010;
        rom[50][5] = 16'h0011;
        rom[50][6] = 16'h003A;
        rom[50][7] = 16'h0019;
        rom[50][8] = 16'h000B;
        rom[50][9] = 16'hFF98;
        rom[50][10] = 16'hFFEA;
        rom[50][11] = 16'h000C;
        rom[50][12] = 16'h001C;
        rom[50][13] = 16'h0019;
        rom[50][14] = 16'hFFBF;
        rom[50][15] = 16'hFFCE;
        rom[50][16] = 16'h002D;
        rom[50][17] = 16'h003C;
        rom[50][18] = 16'hFFCD;
        rom[50][19] = 16'h0033;
        rom[50][20] = 16'hFFD6;
        rom[50][21] = 16'hFFFB;
        rom[50][22] = 16'h0038;
        rom[50][23] = 16'h0011;
        rom[50][24] = 16'hFFC4;
        rom[50][25] = 16'hFFE4;
        rom[50][26] = 16'h0019;
        rom[50][27] = 16'hFFF0;
        rom[50][28] = 16'hFFEF;
        rom[50][29] = 16'hFFE2;
        rom[50][30] = 16'hFFFA;
        rom[50][31] = 16'hFFE8;
        rom[50][32] = 16'hFFFE;
        rom[50][33] = 16'hFFD8;
        rom[50][34] = 16'hFFF9;
        rom[50][35] = 16'hFFEF;
        rom[50][36] = 16'h0029;
        rom[50][37] = 16'h0032;
        rom[50][38] = 16'hFFBF;
        rom[50][39] = 16'hFFF8;
        rom[50][40] = 16'hFFCD;
        rom[50][41] = 16'hFFE9;
        rom[50][42] = 16'h0015;
        rom[50][43] = 16'hFFE7;
        rom[50][44] = 16'h0014;
        rom[50][45] = 16'h0020;
        rom[50][46] = 16'hFFF7;
        rom[50][47] = 16'hFFB9;
        rom[50][48] = 16'h0046;
        rom[50][49] = 16'hFFEE;
        rom[50][50] = 16'hFFF8;
        rom[50][51] = 16'hFFEA;
        rom[50][52] = 16'h0009;
        rom[50][53] = 16'h0032;
        rom[50][54] = 16'hFFCB;
        rom[50][55] = 16'hFFE0;
        rom[50][56] = 16'h0003;
        rom[50][57] = 16'h0003;
        rom[50][58] = 16'hFFF1;
        rom[50][59] = 16'h0002;
        rom[50][60] = 16'h0011;
        rom[50][61] = 16'hFFE1;
        rom[50][62] = 16'hFFFF;
        rom[50][63] = 16'hFFE8;
        rom[50][64] = 16'hFFBC;
        rom[50][65] = 16'hFFE6;
        rom[50][66] = 16'h0011;
        rom[50][67] = 16'hFFF7;
        rom[50][68] = 16'h0013;
        rom[50][69] = 16'hFFF7;
        rom[50][70] = 16'hFFD2;
        rom[50][71] = 16'h0021;
        rom[50][72] = 16'h000F;
        rom[50][73] = 16'hFFDB;
        rom[50][74] = 16'hFFF0;
        rom[50][75] = 16'hFFD5;
        rom[50][76] = 16'h001A;
        rom[50][77] = 16'h0001;
        rom[50][78] = 16'hFFE4;
        rom[50][79] = 16'hFFDF;
        rom[50][80] = 16'hFFEF;
        rom[50][81] = 16'hFFFE;
        rom[50][82] = 16'h0025;
        rom[50][83] = 16'hFFC4;
        rom[50][84] = 16'hFFCF;
        rom[50][85] = 16'hFFC5;
        rom[50][86] = 16'hFFC5;
        rom[50][87] = 16'h0002;
        rom[50][88] = 16'hFFD2;
        rom[50][89] = 16'hFFD4;
        rom[50][90] = 16'h0028;
        rom[50][91] = 16'h004A;
        rom[50][92] = 16'h0022;
        rom[50][93] = 16'h000B;
        rom[50][94] = 16'hFFFF;
        rom[50][95] = 16'hFFEC;
        rom[50][96] = 16'h0004;
        rom[50][97] = 16'h001F;
        rom[50][98] = 16'hFFFA;
        rom[50][99] = 16'h0024;
        rom[50][100] = 16'h0031;
        rom[50][101] = 16'hFFE4;
        rom[50][102] = 16'h0011;
        rom[50][103] = 16'h001C;
        rom[50][104] = 16'h0011;
        rom[50][105] = 16'h000D;
        rom[50][106] = 16'h0006;
        rom[50][107] = 16'hFFF6;
        rom[50][108] = 16'h0017;
        rom[50][109] = 16'hFFE9;
        rom[50][110] = 16'h0006;
        rom[50][111] = 16'h001A;
        rom[50][112] = 16'hFFBD;
        rom[50][113] = 16'h0007;
        rom[50][114] = 16'h0030;
        rom[50][115] = 16'h001C;
        rom[50][116] = 16'h0011;
        rom[50][117] = 16'h0003;
        rom[50][118] = 16'hFFF4;
        rom[50][119] = 16'hFFF5;
        rom[50][120] = 16'hFFEE;
        rom[50][121] = 16'hFFF7;
        rom[50][122] = 16'h0016;
        rom[50][123] = 16'hFFE6;
        rom[50][124] = 16'hFFF9;
        rom[50][125] = 16'hFFE0;
        rom[50][126] = 16'hFFF2;
        rom[50][127] = 16'h001F;
        rom[51][0] = 16'hFFFA;
        rom[51][1] = 16'hFFD4;
        rom[51][2] = 16'h0012;
        rom[51][3] = 16'hFFF5;
        rom[51][4] = 16'h0017;
        rom[51][5] = 16'h000C;
        rom[51][6] = 16'h000D;
        rom[51][7] = 16'hFFC5;
        rom[51][8] = 16'hFFEF;
        rom[51][9] = 16'h002C;
        rom[51][10] = 16'h0000;
        rom[51][11] = 16'h002A;
        rom[51][12] = 16'hFFD4;
        rom[51][13] = 16'hFFE9;
        rom[51][14] = 16'hFFFF;
        rom[51][15] = 16'h0031;
        rom[51][16] = 16'h0033;
        rom[51][17] = 16'hFFE2;
        rom[51][18] = 16'h000D;
        rom[51][19] = 16'hFFD8;
        rom[51][20] = 16'hFFE8;
        rom[51][21] = 16'h001F;
        rom[51][22] = 16'h000D;
        rom[51][23] = 16'h000D;
        rom[51][24] = 16'h001F;
        rom[51][25] = 16'hFFEE;
        rom[51][26] = 16'hFFE5;
        rom[51][27] = 16'hFFEA;
        rom[51][28] = 16'hFFD2;
        rom[51][29] = 16'hFFEF;
        rom[51][30] = 16'hFFFE;
        rom[51][31] = 16'h0007;
        rom[51][32] = 16'h0005;
        rom[51][33] = 16'hFFFE;
        rom[51][34] = 16'h0024;
        rom[51][35] = 16'hFFF4;
        rom[51][36] = 16'hFFD3;
        rom[51][37] = 16'hFFEF;
        rom[51][38] = 16'h0011;
        rom[51][39] = 16'hFFEB;
        rom[51][40] = 16'hFFE2;
        rom[51][41] = 16'h0002;
        rom[51][42] = 16'hFFF6;
        rom[51][43] = 16'h0014;
        rom[51][44] = 16'hFFB0;
        rom[51][45] = 16'hFFD8;
        rom[51][46] = 16'h0011;
        rom[51][47] = 16'h0013;
        rom[51][48] = 16'hFFC8;
        rom[51][49] = 16'hFFE9;
        rom[51][50] = 16'h001A;
        rom[51][51] = 16'hFFFD;
        rom[51][52] = 16'h000E;
        rom[51][53] = 16'hFFE4;
        rom[51][54] = 16'h0009;
        rom[51][55] = 16'hFFFD;
        rom[51][56] = 16'h0013;
        rom[51][57] = 16'hFFE1;
        rom[51][58] = 16'hFFFF;
        rom[51][59] = 16'hFFFE;
        rom[51][60] = 16'hFFF9;
        rom[51][61] = 16'hFFEC;
        rom[51][62] = 16'hFFF6;
        rom[51][63] = 16'hFFC0;
        rom[51][64] = 16'hFFF9;
        rom[51][65] = 16'hFFE5;
        rom[51][66] = 16'hFFF3;
        rom[51][67] = 16'hFFFE;
        rom[51][68] = 16'hFFD1;
        rom[51][69] = 16'hFFE6;
        rom[51][70] = 16'h000D;
        rom[51][71] = 16'hFFF4;
        rom[51][72] = 16'h0016;
        rom[51][73] = 16'h0007;
        rom[51][74] = 16'hFFDF;
        rom[51][75] = 16'h0018;
        rom[51][76] = 16'h0015;
        rom[51][77] = 16'hFFF9;
        rom[51][78] = 16'hFFB5;
        rom[51][79] = 16'h0016;
        rom[51][80] = 16'hFFB6;
        rom[51][81] = 16'hFFFE;
        rom[51][82] = 16'hFFF9;
        rom[51][83] = 16'h0016;
        rom[51][84] = 16'hFFEF;
        rom[51][85] = 16'hFFA4;
        rom[51][86] = 16'h0007;
        rom[51][87] = 16'h0017;
        rom[51][88] = 16'hFFC5;
        rom[51][89] = 16'hFFD4;
        rom[51][90] = 16'h0003;
        rom[51][91] = 16'hFFEF;
        rom[51][92] = 16'h0033;
        rom[51][93] = 16'hFFBE;
        rom[51][94] = 16'hFFDB;
        rom[51][95] = 16'hFFED;
        rom[51][96] = 16'h001B;
        rom[51][97] = 16'h0033;
        rom[51][98] = 16'hFFE8;
        rom[51][99] = 16'hFFF5;
        rom[51][100] = 16'h0002;
        rom[51][101] = 16'hFFEE;
        rom[51][102] = 16'h0019;
        rom[51][103] = 16'h000D;
        rom[51][104] = 16'hFFCF;
        rom[51][105] = 16'h0016;
        rom[51][106] = 16'hFFFF;
        rom[51][107] = 16'hFFF8;
        rom[51][108] = 16'h002C;
        rom[51][109] = 16'hFFEC;
        rom[51][110] = 16'h001D;
        rom[51][111] = 16'hFFC7;
        rom[51][112] = 16'hFFE5;
        rom[51][113] = 16'hFFFD;
        rom[51][114] = 16'h0021;
        rom[51][115] = 16'hFFEA;
        rom[51][116] = 16'h000F;
        rom[51][117] = 16'hFFFB;
        rom[51][118] = 16'hFFE8;
        rom[51][119] = 16'h0004;
        rom[51][120] = 16'h0031;
        rom[51][121] = 16'h001F;
        rom[51][122] = 16'h002C;
        rom[51][123] = 16'h0018;
        rom[51][124] = 16'h0007;
        rom[51][125] = 16'h001F;
        rom[51][126] = 16'hFFDF;
        rom[51][127] = 16'hFFE8;
        rom[52][0] = 16'hFFFE;
        rom[52][1] = 16'hFFDE;
        rom[52][2] = 16'hFFB0;
        rom[52][3] = 16'h001B;
        rom[52][4] = 16'hFFB9;
        rom[52][5] = 16'hFFCF;
        rom[52][6] = 16'hFFDE;
        rom[52][7] = 16'h0002;
        rom[52][8] = 16'h0002;
        rom[52][9] = 16'hFFD8;
        rom[52][10] = 16'hFFF8;
        rom[52][11] = 16'h0013;
        rom[52][12] = 16'h0019;
        rom[52][13] = 16'h001C;
        rom[52][14] = 16'hFFCD;
        rom[52][15] = 16'h0011;
        rom[52][16] = 16'hFFF1;
        rom[52][17] = 16'h0006;
        rom[52][18] = 16'hFFD3;
        rom[52][19] = 16'hFFE5;
        rom[52][20] = 16'hFFE7;
        rom[52][21] = 16'h001C;
        rom[52][22] = 16'h0000;
        rom[52][23] = 16'h001A;
        rom[52][24] = 16'h0020;
        rom[52][25] = 16'hFFED;
        rom[52][26] = 16'hFFEB;
        rom[52][27] = 16'hFFFC;
        rom[52][28] = 16'h000E;
        rom[52][29] = 16'h0010;
        rom[52][30] = 16'hFFF4;
        rom[52][31] = 16'hFFEF;
        rom[52][32] = 16'hFFA9;
        rom[52][33] = 16'hFFF3;
        rom[52][34] = 16'h0000;
        rom[52][35] = 16'h002F;
        rom[52][36] = 16'hFFC2;
        rom[52][37] = 16'h0014;
        rom[52][38] = 16'hFFB7;
        rom[52][39] = 16'h001F;
        rom[52][40] = 16'h000D;
        rom[52][41] = 16'h0016;
        rom[52][42] = 16'h0025;
        rom[52][43] = 16'hFFF6;
        rom[52][44] = 16'h0010;
        rom[52][45] = 16'h0009;
        rom[52][46] = 16'h0002;
        rom[52][47] = 16'h0021;
        rom[52][48] = 16'hFFF9;
        rom[52][49] = 16'hFFE1;
        rom[52][50] = 16'hFFD2;
        rom[52][51] = 16'hFFF9;
        rom[52][52] = 16'hFFC3;
        rom[52][53] = 16'hFFDF;
        rom[52][54] = 16'hFFDC;
        rom[52][55] = 16'h0024;
        rom[52][56] = 16'hFFFE;
        rom[52][57] = 16'hFFFA;
        rom[52][58] = 16'h001F;
        rom[52][59] = 16'h000C;
        rom[52][60] = 16'hFFE2;
        rom[52][61] = 16'h0004;
        rom[52][62] = 16'hFFDC;
        rom[52][63] = 16'h000A;
        rom[52][64] = 16'h000F;
        rom[52][65] = 16'hFFEF;
        rom[52][66] = 16'hFFCB;
        rom[52][67] = 16'hFFD5;
        rom[52][68] = 16'h000B;
        rom[52][69] = 16'h0011;
        rom[52][70] = 16'hFFC8;
        rom[52][71] = 16'hFFE0;
        rom[52][72] = 16'hFFF2;
        rom[52][73] = 16'hFFF1;
        rom[52][74] = 16'h0021;
        rom[52][75] = 16'hFFF6;
        rom[52][76] = 16'h0003;
        rom[52][77] = 16'h001F;
        rom[52][78] = 16'h0011;
        rom[52][79] = 16'hFFE4;
        rom[52][80] = 16'h000E;
        rom[52][81] = 16'hFFF0;
        rom[52][82] = 16'hFFFA;
        rom[52][83] = 16'h0033;
        rom[52][84] = 16'hFFF2;
        rom[52][85] = 16'hFFC2;
        rom[52][86] = 16'h0007;
        rom[52][87] = 16'hFFDC;
        rom[52][88] = 16'hFFE4;
        rom[52][89] = 16'hFFEB;
        rom[52][90] = 16'hFFDF;
        rom[52][91] = 16'h0003;
        rom[52][92] = 16'h0032;
        rom[52][93] = 16'h0011;
        rom[52][94] = 16'h000A;
        rom[52][95] = 16'hFFFE;
        rom[52][96] = 16'hFFE3;
        rom[52][97] = 16'hFFD7;
        rom[52][98] = 16'h0001;
        rom[52][99] = 16'h0008;
        rom[52][100] = 16'h0016;
        rom[52][101] = 16'hFFEE;
        rom[52][102] = 16'h0009;
        rom[52][103] = 16'h0026;
        rom[52][104] = 16'hFFF4;
        rom[52][105] = 16'hFFF4;
        rom[52][106] = 16'hFFF9;
        rom[52][107] = 16'hFFE1;
        rom[52][108] = 16'hFFCD;
        rom[52][109] = 16'h0016;
        rom[52][110] = 16'hFFFE;
        rom[52][111] = 16'h001B;
        rom[52][112] = 16'h0018;
        rom[52][113] = 16'h002D;
        rom[52][114] = 16'hFFFD;
        rom[52][115] = 16'hFFCE;
        rom[52][116] = 16'hFFF1;
        rom[52][117] = 16'hFFE2;
        rom[52][118] = 16'h0005;
        rom[52][119] = 16'hFFDA;
        rom[52][120] = 16'h0000;
        rom[52][121] = 16'hFFF4;
        rom[52][122] = 16'h0025;
        rom[52][123] = 16'h0014;
        rom[52][124] = 16'hFFD7;
        rom[52][125] = 16'hFFFF;
        rom[52][126] = 16'hFFF9;
        rom[52][127] = 16'hFFEF;
        rom[53][0] = 16'hFFE9;
        rom[53][1] = 16'h0011;
        rom[53][2] = 16'hFFF7;
        rom[53][3] = 16'hFFE4;
        rom[53][4] = 16'h0002;
        rom[53][5] = 16'h0021;
        rom[53][6] = 16'h0011;
        rom[53][7] = 16'h0018;
        rom[53][8] = 16'hFFE4;
        rom[53][9] = 16'hFFE3;
        rom[53][10] = 16'hFFF5;
        rom[53][11] = 16'hFFE7;
        rom[53][12] = 16'hFFE7;
        rom[53][13] = 16'hFFE8;
        rom[53][14] = 16'h0006;
        rom[53][15] = 16'hFFF4;
        rom[53][16] = 16'hFFFD;
        rom[53][17] = 16'h0004;
        rom[53][18] = 16'hFFE3;
        rom[53][19] = 16'hFFDA;
        rom[53][20] = 16'hFFFB;
        rom[53][21] = 16'hFFF4;
        rom[53][22] = 16'h000B;
        rom[53][23] = 16'hFFE7;
        rom[53][24] = 16'h0006;
        rom[53][25] = 16'hFFEA;
        rom[53][26] = 16'h0012;
        rom[53][27] = 16'hFFCB;
        rom[53][28] = 16'h001D;
        rom[53][29] = 16'hFFF7;
        rom[53][30] = 16'hFFCD;
        rom[53][31] = 16'hFFEF;
        rom[53][32] = 16'h000F;
        rom[53][33] = 16'h000E;
        rom[53][34] = 16'hFFC0;
        rom[53][35] = 16'h002C;
        rom[53][36] = 16'h0015;
        rom[53][37] = 16'hFFF9;
        rom[53][38] = 16'h0008;
        rom[53][39] = 16'hFFD2;
        rom[53][40] = 16'hFFEA;
        rom[53][41] = 16'hFFE0;
        rom[53][42] = 16'h0009;
        rom[53][43] = 16'h0003;
        rom[53][44] = 16'hFFEA;
        rom[53][45] = 16'h001F;
        rom[53][46] = 16'h000C;
        rom[53][47] = 16'h0009;
        rom[53][48] = 16'h0002;
        rom[53][49] = 16'hFFF6;
        rom[53][50] = 16'h0025;
        rom[53][51] = 16'hFFC1;
        rom[53][52] = 16'hFFEA;
        rom[53][53] = 16'hFFB5;
        rom[53][54] = 16'h0032;
        rom[53][55] = 16'hFFEF;
        rom[53][56] = 16'hFFF0;
        rom[53][57] = 16'hFFB3;
        rom[53][58] = 16'h0016;
        rom[53][59] = 16'hFFE4;
        rom[53][60] = 16'hFFEA;
        rom[53][61] = 16'h0019;
        rom[53][62] = 16'h0033;
        rom[53][63] = 16'h0006;
        rom[53][64] = 16'hFFED;
        rom[53][65] = 16'h0014;
        rom[53][66] = 16'hFFF3;
        rom[53][67] = 16'hFFEE;
        rom[53][68] = 16'hFFE7;
        rom[53][69] = 16'hFFE7;
        rom[53][70] = 16'hFFFA;
        rom[53][71] = 16'h0025;
        rom[53][72] = 16'hFFF4;
        rom[53][73] = 16'hFFEF;
        rom[53][74] = 16'h0006;
        rom[53][75] = 16'h0018;
        rom[53][76] = 16'hFFDD;
        rom[53][77] = 16'h0059;
        rom[53][78] = 16'hFFFF;
        rom[53][79] = 16'hFFF4;
        rom[53][80] = 16'h000C;
        rom[53][81] = 16'h0018;
        rom[53][82] = 16'h0016;
        rom[53][83] = 16'h000B;
        rom[53][84] = 16'h0004;
        rom[53][85] = 16'hFFEA;
        rom[53][86] = 16'hFFCF;
        rom[53][87] = 16'hFFCC;
        rom[53][88] = 16'hFFDE;
        rom[53][89] = 16'h0002;
        rom[53][90] = 16'hFFF1;
        rom[53][91] = 16'h0016;
        rom[53][92] = 16'hFFFD;
        rom[53][93] = 16'h0018;
        rom[53][94] = 16'hFFEF;
        rom[53][95] = 16'hFFDA;
        rom[53][96] = 16'h0012;
        rom[53][97] = 16'hFFF7;
        rom[53][98] = 16'hFFF2;
        rom[53][99] = 16'h0011;
        rom[53][100] = 16'h0033;
        rom[53][101] = 16'h0023;
        rom[53][102] = 16'h0022;
        rom[53][103] = 16'hFFF7;
        rom[53][104] = 16'hFF96;
        rom[53][105] = 16'hFFD7;
        rom[53][106] = 16'hFFE8;
        rom[53][107] = 16'h0011;
        rom[53][108] = 16'h0023;
        rom[53][109] = 16'h0046;
        rom[53][110] = 16'h000C;
        rom[53][111] = 16'h000A;
        rom[53][112] = 16'h000C;
        rom[53][113] = 16'hFFF8;
        rom[53][114] = 16'h0013;
        rom[53][115] = 16'hFFE6;
        rom[53][116] = 16'h0033;
        rom[53][117] = 16'hFFD0;
        rom[53][118] = 16'h000C;
        rom[53][119] = 16'h0017;
        rom[53][120] = 16'hFFC5;
        rom[53][121] = 16'hFFDC;
        rom[53][122] = 16'hFFC8;
        rom[53][123] = 16'hFFEA;
        rom[53][124] = 16'h0001;
        rom[53][125] = 16'hFFBD;
        rom[53][126] = 16'hFFE5;
        rom[53][127] = 16'hFFB7;
        rom[54][0] = 16'h001B;
        rom[54][1] = 16'hFFEB;
        rom[54][2] = 16'hFFF5;
        rom[54][3] = 16'hFFB5;
        rom[54][4] = 16'hFFE1;
        rom[54][5] = 16'hFFD2;
        rom[54][6] = 16'hFFB0;
        rom[54][7] = 16'hFFFB;
        rom[54][8] = 16'h0016;
        rom[54][9] = 16'hFFE8;
        rom[54][10] = 16'hFFE1;
        rom[54][11] = 16'h0002;
        rom[54][12] = 16'h0022;
        rom[54][13] = 16'h001C;
        rom[54][14] = 16'hFFD0;
        rom[54][15] = 16'hFFF6;
        rom[54][16] = 16'h0007;
        rom[54][17] = 16'h0022;
        rom[54][18] = 16'h0003;
        rom[54][19] = 16'h0003;
        rom[54][20] = 16'hFFF5;
        rom[54][21] = 16'hFFF3;
        rom[54][22] = 16'h0002;
        rom[54][23] = 16'h000C;
        rom[54][24] = 16'h0003;
        rom[54][25] = 16'hFFCA;
        rom[54][26] = 16'hFFBC;
        rom[54][27] = 16'h001C;
        rom[54][28] = 16'hFFD7;
        rom[54][29] = 16'hFFF8;
        rom[54][30] = 16'h0007;
        rom[54][31] = 16'hFFEF;
        rom[54][32] = 16'h0002;
        rom[54][33] = 16'h0010;
        rom[54][34] = 16'hFFFA;
        rom[54][35] = 16'hFFFB;
        rom[54][36] = 16'hFFF3;
        rom[54][37] = 16'hFFE5;
        rom[54][38] = 16'h001E;
        rom[54][39] = 16'h0002;
        rom[54][40] = 16'hFFE7;
        rom[54][41] = 16'hFFF3;
        rom[54][42] = 16'h002A;
        rom[54][43] = 16'hFFDC;
        rom[54][44] = 16'h002F;
        rom[54][45] = 16'h0012;
        rom[54][46] = 16'hFFFD;
        rom[54][47] = 16'hFFEB;
        rom[54][48] = 16'hFFFA;
        rom[54][49] = 16'hFFEE;
        rom[54][50] = 16'h0017;
        rom[54][51] = 16'h000A;
        rom[54][52] = 16'hFFF1;
        rom[54][53] = 16'hFFF7;
        rom[54][54] = 16'hFFE7;
        rom[54][55] = 16'hFFB7;
        rom[54][56] = 16'h0029;
        rom[54][57] = 16'h0018;
        rom[54][58] = 16'h0016;
        rom[54][59] = 16'hFFFD;
        rom[54][60] = 16'hFFF1;
        rom[54][61] = 16'hFFF9;
        rom[54][62] = 16'hFFEC;
        rom[54][63] = 16'hFFD2;
        rom[54][64] = 16'hFFB0;
        rom[54][65] = 16'h0007;
        rom[54][66] = 16'hFFCA;
        rom[54][67] = 16'hFFCB;
        rom[54][68] = 16'hFFC5;
        rom[54][69] = 16'hFFDA;
        rom[54][70] = 16'h0016;
        rom[54][71] = 16'hFFC8;
        rom[54][72] = 16'h0007;
        rom[54][73] = 16'hFFEC;
        rom[54][74] = 16'h0002;
        rom[54][75] = 16'h0010;
        rom[54][76] = 16'h0019;
        rom[54][77] = 16'h0015;
        rom[54][78] = 16'hFFFC;
        rom[54][79] = 16'hFFFE;
        rom[54][80] = 16'hFFDA;
        rom[54][81] = 16'h002B;
        rom[54][82] = 16'hFFBA;
        rom[54][83] = 16'h002E;
        rom[54][84] = 16'hFFFC;
        rom[54][85] = 16'h0008;
        rom[54][86] = 16'hFFF6;
        rom[54][87] = 16'hFFE2;
        rom[54][88] = 16'hFFEF;
        rom[54][89] = 16'h0026;
        rom[54][90] = 16'hFFE2;
        rom[54][91] = 16'h0002;
        rom[54][92] = 16'hFFFD;
        rom[54][93] = 16'h0001;
        rom[54][94] = 16'h000E;
        rom[54][95] = 16'hFFEB;
        rom[54][96] = 16'hFFB9;
        rom[54][97] = 16'hFFBB;
        rom[54][98] = 16'hFFFA;
        rom[54][99] = 16'h0011;
        rom[54][100] = 16'hFFB3;
        rom[54][101] = 16'hFFCE;
        rom[54][102] = 16'hFFEB;
        rom[54][103] = 16'hFFE1;
        rom[54][104] = 16'hFFD4;
        rom[54][105] = 16'hFFD5;
        rom[54][106] = 16'hFFED;
        rom[54][107] = 16'h000D;
        rom[54][108] = 16'h0007;
        rom[54][109] = 16'hFFDD;
        rom[54][110] = 16'h000D;
        rom[54][111] = 16'h0008;
        rom[54][112] = 16'h0042;
        rom[54][113] = 16'h0002;
        rom[54][114] = 16'h0002;
        rom[54][115] = 16'hFFC6;
        rom[54][116] = 16'hFFF2;
        rom[54][117] = 16'hFFAE;
        rom[54][118] = 16'hFFFA;
        rom[54][119] = 16'hFFFF;
        rom[54][120] = 16'hFFFA;
        rom[54][121] = 16'hFFC4;
        rom[54][122] = 16'h0013;
        rom[54][123] = 16'h001E;
        rom[54][124] = 16'hFFFE;
        rom[54][125] = 16'hFFF2;
        rom[54][126] = 16'hFFE2;
        rom[54][127] = 16'hFFFC;
        rom[55][0] = 16'h000B;
        rom[55][1] = 16'h0003;
        rom[55][2] = 16'hFFD7;
        rom[55][3] = 16'hFFD9;
        rom[55][4] = 16'h0010;
        rom[55][5] = 16'hFFE4;
        rom[55][6] = 16'h0011;
        rom[55][7] = 16'h0018;
        rom[55][8] = 16'h001B;
        rom[55][9] = 16'hFFF7;
        rom[55][10] = 16'h001F;
        rom[55][11] = 16'h0015;
        rom[55][12] = 16'hFFE1;
        rom[55][13] = 16'hFFDD;
        rom[55][14] = 16'h0026;
        rom[55][15] = 16'hFFF4;
        rom[55][16] = 16'hFFC8;
        rom[55][17] = 16'h0029;
        rom[55][18] = 16'h001E;
        rom[55][19] = 16'h0003;
        rom[55][20] = 16'hFFFE;
        rom[55][21] = 16'hFFF0;
        rom[55][22] = 16'h0005;
        rom[55][23] = 16'h0002;
        rom[55][24] = 16'hFFE0;
        rom[55][25] = 16'hFFCD;
        rom[55][26] = 16'h0027;
        rom[55][27] = 16'hFFE1;
        rom[55][28] = 16'hFFF3;
        rom[55][29] = 16'hFFFE;
        rom[55][30] = 16'h000C;
        rom[55][31] = 16'hFFF1;
        rom[55][32] = 16'hFFFF;
        rom[55][33] = 16'h0028;
        rom[55][34] = 16'hFFEC;
        rom[55][35] = 16'h0002;
        rom[55][36] = 16'hFFAD;
        rom[55][37] = 16'hFFED;
        rom[55][38] = 16'hFFFF;
        rom[55][39] = 16'h0016;
        rom[55][40] = 16'hFFDB;
        rom[55][41] = 16'h001B;
        rom[55][42] = 16'hFFFE;
        rom[55][43] = 16'h0018;
        rom[55][44] = 16'hFFDC;
        rom[55][45] = 16'h0009;
        rom[55][46] = 16'hFFBF;
        rom[55][47] = 16'hFFB1;
        rom[55][48] = 16'hFFCA;
        rom[55][49] = 16'hFFD4;
        rom[55][50] = 16'hFFB7;
        rom[55][51] = 16'h0014;
        rom[55][52] = 16'hFFFB;
        rom[55][53] = 16'h001C;
        rom[55][54] = 16'hFFFB;
        rom[55][55] = 16'hFFDC;
        rom[55][56] = 16'hFFE1;
        rom[55][57] = 16'h0012;
        rom[55][58] = 16'h0002;
        rom[55][59] = 16'h000D;
        rom[55][60] = 16'hFFD5;
        rom[55][61] = 16'h0003;
        rom[55][62] = 16'hFFFC;
        rom[55][63] = 16'h001E;
        rom[55][64] = 16'hFFDE;
        rom[55][65] = 16'hFFDB;
        rom[55][66] = 16'hFFF4;
        rom[55][67] = 16'h0006;
        rom[55][68] = 16'h0046;
        rom[55][69] = 16'hFFD8;
        rom[55][70] = 16'h000B;
        rom[55][71] = 16'h0024;
        rom[55][72] = 16'h000C;
        rom[55][73] = 16'hFFEF;
        rom[55][74] = 16'h000E;
        rom[55][75] = 16'h0026;
        rom[55][76] = 16'hFFE8;
        rom[55][77] = 16'h001B;
        rom[55][78] = 16'hFFF1;
        rom[55][79] = 16'hFFD7;
        rom[55][80] = 16'hFFE8;
        rom[55][81] = 16'h000B;
        rom[55][82] = 16'hFFD8;
        rom[55][83] = 16'hFFFC;
        rom[55][84] = 16'hFFC5;
        rom[55][85] = 16'hFFB4;
        rom[55][86] = 16'h0012;
        rom[55][87] = 16'hFFFA;
        rom[55][88] = 16'hFFD2;
        rom[55][89] = 16'h001F;
        rom[55][90] = 16'hFFE6;
        rom[55][91] = 16'hFFDE;
        rom[55][92] = 16'hFFD8;
        rom[55][93] = 16'h001B;
        rom[55][94] = 16'h0004;
        rom[55][95] = 16'h000C;
        rom[55][96] = 16'h0026;
        rom[55][97] = 16'h0029;
        rom[55][98] = 16'hFFC8;
        rom[55][99] = 16'hFFFF;
        rom[55][100] = 16'h000C;
        rom[55][101] = 16'h0029;
        rom[55][102] = 16'hFFE3;
        rom[55][103] = 16'h0013;
        rom[55][104] = 16'hFFF8;
        rom[55][105] = 16'h0001;
        rom[55][106] = 16'hFFC1;
        rom[55][107] = 16'h0019;
        rom[55][108] = 16'hFFEA;
        rom[55][109] = 16'hFFFE;
        rom[55][110] = 16'hFFD1;
        rom[55][111] = 16'hFFDB;
        rom[55][112] = 16'h001F;
        rom[55][113] = 16'hFFE3;
        rom[55][114] = 16'hFFEF;
        rom[55][115] = 16'hFFD9;
        rom[55][116] = 16'h0002;
        rom[55][117] = 16'h001E;
        rom[55][118] = 16'hFFF9;
        rom[55][119] = 16'hFFEB;
        rom[55][120] = 16'hFFE4;
        rom[55][121] = 16'hFFEF;
        rom[55][122] = 16'h000D;
        rom[55][123] = 16'hFFA5;
        rom[55][124] = 16'h0002;
        rom[55][125] = 16'hFFE4;
        rom[55][126] = 16'h001B;
        rom[55][127] = 16'h0014;
        rom[56][0] = 16'h0022;
        rom[56][1] = 16'h0007;
        rom[56][2] = 16'hFFF8;
        rom[56][3] = 16'hFFDE;
        rom[56][4] = 16'hFFFE;
        rom[56][5] = 16'h0016;
        rom[56][6] = 16'h0002;
        rom[56][7] = 16'h0012;
        rom[56][8] = 16'h0011;
        rom[56][9] = 16'hFFFC;
        rom[56][10] = 16'hFFF9;
        rom[56][11] = 16'hFFBA;
        rom[56][12] = 16'hFFD9;
        rom[56][13] = 16'hFFE9;
        rom[56][14] = 16'hFFF5;
        rom[56][15] = 16'h001E;
        rom[56][16] = 16'hFFF9;
        rom[56][17] = 16'hFFAB;
        rom[56][18] = 16'hFFDF;
        rom[56][19] = 16'h0027;
        rom[56][20] = 16'hFFEB;
        rom[56][21] = 16'hFFF3;
        rom[56][22] = 16'hFFD1;
        rom[56][23] = 16'hFFE3;
        rom[56][24] = 16'h004B;
        rom[56][25] = 16'h0001;
        rom[56][26] = 16'hFFEF;
        rom[56][27] = 16'hFFC9;
        rom[56][28] = 16'h000F;
        rom[56][29] = 16'h0001;
        rom[56][30] = 16'hFFE5;
        rom[56][31] = 16'hFFFE;
        rom[56][32] = 16'h0013;
        rom[56][33] = 16'h002C;
        rom[56][34] = 16'h0002;
        rom[56][35] = 16'h0008;
        rom[56][36] = 16'hFFFE;
        rom[56][37] = 16'hFFF9;
        rom[56][38] = 16'h004C;
        rom[56][39] = 16'h0018;
        rom[56][40] = 16'hFFDA;
        rom[56][41] = 16'h0002;
        rom[56][42] = 16'hFFDD;
        rom[56][43] = 16'hFFC3;
        rom[56][44] = 16'h0017;
        rom[56][45] = 16'h000E;
        rom[56][46] = 16'hFFF3;
        rom[56][47] = 16'hFFFE;
        rom[56][48] = 16'h0016;
        rom[56][49] = 16'h001E;
        rom[56][50] = 16'hFFF3;
        rom[56][51] = 16'hFFE5;
        rom[56][52] = 16'hFFF0;
        rom[56][53] = 16'hFFE6;
        rom[56][54] = 16'hFFD8;
        rom[56][55] = 16'hFFF6;
        rom[56][56] = 16'h0000;
        rom[56][57] = 16'h000C;
        rom[56][58] = 16'hFFFE;
        rom[56][59] = 16'hFFC5;
        rom[56][60] = 16'hFFDB;
        rom[56][61] = 16'h0000;
        rom[56][62] = 16'hFFF8;
        rom[56][63] = 16'h001C;
        rom[56][64] = 16'h0006;
        rom[56][65] = 16'hFFF0;
        rom[56][66] = 16'hFFD1;
        rom[56][67] = 16'hFFFD;
        rom[56][68] = 16'hFFD9;
        rom[56][69] = 16'hFFFA;
        rom[56][70] = 16'h000B;
        rom[56][71] = 16'hFFD6;
        rom[56][72] = 16'hFFFF;
        rom[56][73] = 16'hFFF5;
        rom[56][74] = 16'hFFE1;
        rom[56][75] = 16'h003C;
        rom[56][76] = 16'hFFFA;
        rom[56][77] = 16'hFFC1;
        rom[56][78] = 16'h0005;
        rom[56][79] = 16'hFFF9;
        rom[56][80] = 16'hFFD2;
        rom[56][81] = 16'h0000;
        rom[56][82] = 16'h0002;
        rom[56][83] = 16'h0029;
        rom[56][84] = 16'h0004;
        rom[56][85] = 16'hFFEB;
        rom[56][86] = 16'h0019;
        rom[56][87] = 16'hFFBF;
        rom[56][88] = 16'h0000;
        rom[56][89] = 16'hFFDE;
        rom[56][90] = 16'h0009;
        rom[56][91] = 16'hFFFC;
        rom[56][92] = 16'hFFF1;
        rom[56][93] = 16'hFFEE;
        rom[56][94] = 16'hFFB8;
        rom[56][95] = 16'h0010;
        rom[56][96] = 16'hFFDA;
        rom[56][97] = 16'h000D;
        rom[56][98] = 16'hFFEC;
        rom[56][99] = 16'h000B;
        rom[56][100] = 16'h0006;
        rom[56][101] = 16'hFFD3;
        rom[56][102] = 16'h0010;
        rom[56][103] = 16'hFFF9;
        rom[56][104] = 16'hFFD4;
        rom[56][105] = 16'h0019;
        rom[56][106] = 16'hFFE2;
        rom[56][107] = 16'h000C;
        rom[56][108] = 16'h000A;
        rom[56][109] = 16'hFFE1;
        rom[56][110] = 16'h0003;
        rom[56][111] = 16'h0014;
        rom[56][112] = 16'hFFDB;
        rom[56][113] = 16'h0000;
        rom[56][114] = 16'h0002;
        rom[56][115] = 16'hFFF9;
        rom[56][116] = 16'hFFF3;
        rom[56][117] = 16'hFFE8;
        rom[56][118] = 16'hFFFB;
        rom[56][119] = 16'h000E;
        rom[56][120] = 16'hFFEC;
        rom[56][121] = 16'h0003;
        rom[56][122] = 16'hFFBE;
        rom[56][123] = 16'h000A;
        rom[56][124] = 16'hFFDB;
        rom[56][125] = 16'hFFDE;
        rom[56][126] = 16'hFFC0;
        rom[56][127] = 16'h0012;
        rom[57][0] = 16'h0021;
        rom[57][1] = 16'hFFFC;
        rom[57][2] = 16'h0001;
        rom[57][3] = 16'hFFEF;
        rom[57][4] = 16'h0002;
        rom[57][5] = 16'h0005;
        rom[57][6] = 16'hFFCB;
        rom[57][7] = 16'hFFEB;
        rom[57][8] = 16'h0011;
        rom[57][9] = 16'hFFE6;
        rom[57][10] = 16'hFFD1;
        rom[57][11] = 16'h001F;
        rom[57][12] = 16'h0011;
        rom[57][13] = 16'h0024;
        rom[57][14] = 16'hFFE5;
        rom[57][15] = 16'h001A;
        rom[57][16] = 16'h001D;
        rom[57][17] = 16'hFFF6;
        rom[57][18] = 16'h0000;
        rom[57][19] = 16'hFFD0;
        rom[57][20] = 16'h002E;
        rom[57][21] = 16'hFFEE;
        rom[57][22] = 16'hFFE0;
        rom[57][23] = 16'hFFF3;
        rom[57][24] = 16'hFFEE;
        rom[57][25] = 16'hFFD4;
        rom[57][26] = 16'h0018;
        rom[57][27] = 16'hFFE5;
        rom[57][28] = 16'hFFEF;
        rom[57][29] = 16'h0001;
        rom[57][30] = 16'h0016;
        rom[57][31] = 16'hFFC8;
        rom[57][32] = 16'h0007;
        rom[57][33] = 16'hFFF6;
        rom[57][34] = 16'h0018;
        rom[57][35] = 16'hFFE4;
        rom[57][36] = 16'hFFF5;
        rom[57][37] = 16'hFFF5;
        rom[57][38] = 16'hFFCB;
        rom[57][39] = 16'hFFFF;
        rom[57][40] = 16'h0005;
        rom[57][41] = 16'hFFE0;
        rom[57][42] = 16'hFFF4;
        rom[57][43] = 16'hFFFB;
        rom[57][44] = 16'h0011;
        rom[57][45] = 16'hFFE9;
        rom[57][46] = 16'hFFF0;
        rom[57][47] = 16'hFFE8;
        rom[57][48] = 16'hFFF4;
        rom[57][49] = 16'h0007;
        rom[57][50] = 16'h0011;
        rom[57][51] = 16'h0023;
        rom[57][52] = 16'h0016;
        rom[57][53] = 16'h0009;
        rom[57][54] = 16'h0007;
        rom[57][55] = 16'hFFC6;
        rom[57][56] = 16'h001D;
        rom[57][57] = 16'h000B;
        rom[57][58] = 16'hFFFC;
        rom[57][59] = 16'hFFF2;
        rom[57][60] = 16'h0007;
        rom[57][61] = 16'hFFE8;
        rom[57][62] = 16'hFFB9;
        rom[57][63] = 16'hFFD1;
        rom[57][64] = 16'hFFD8;
        rom[57][65] = 16'h0007;
        rom[57][66] = 16'h0015;
        rom[57][67] = 16'hFFF3;
        rom[57][68] = 16'hFFBE;
        rom[57][69] = 16'hFFDB;
        rom[57][70] = 16'hFFF2;
        rom[57][71] = 16'hFFFA;
        rom[57][72] = 16'h000D;
        rom[57][73] = 16'hFFEA;
        rom[57][74] = 16'hFFA8;
        rom[57][75] = 16'hFFD5;
        rom[57][76] = 16'h000D;
        rom[57][77] = 16'hFFE5;
        rom[57][78] = 16'h0025;
        rom[57][79] = 16'h0017;
        rom[57][80] = 16'h0001;
        rom[57][81] = 16'h001D;
        rom[57][82] = 16'h0020;
        rom[57][83] = 16'h0001;
        rom[57][84] = 16'h0003;
        rom[57][85] = 16'h0003;
        rom[57][86] = 16'h000B;
        rom[57][87] = 16'h0024;
        rom[57][88] = 16'hFFE5;
        rom[57][89] = 16'h000F;
        rom[57][90] = 16'hFFFA;
        rom[57][91] = 16'hFFFD;
        rom[57][92] = 16'h0000;
        rom[57][93] = 16'hFFEF;
        rom[57][94] = 16'h0017;
        rom[57][95] = 16'hFFFD;
        rom[57][96] = 16'hFFEA;
        rom[57][97] = 16'hFFF3;
        rom[57][98] = 16'hFFDC;
        rom[57][99] = 16'hFFFA;
        rom[57][100] = 16'hFFBB;
        rom[57][101] = 16'hFFDF;
        rom[57][102] = 16'hFFDC;
        rom[57][103] = 16'hFFE6;
        rom[57][104] = 16'h0009;
        rom[57][105] = 16'hFFC0;
        rom[57][106] = 16'h000B;
        rom[57][107] = 16'h0005;
        rom[57][108] = 16'hFFE7;
        rom[57][109] = 16'hFFE4;
        rom[57][110] = 16'hFFF7;
        rom[57][111] = 16'h0011;
        rom[57][112] = 16'h0008;
        rom[57][113] = 16'hFFF0;
        rom[57][114] = 16'hFFDA;
        rom[57][115] = 16'hFFF5;
        rom[57][116] = 16'h0020;
        rom[57][117] = 16'hFFD6;
        rom[57][118] = 16'hFFE9;
        rom[57][119] = 16'hFFFB;
        rom[57][120] = 16'h002A;
        rom[57][121] = 16'hFFD0;
        rom[57][122] = 16'h0014;
        rom[57][123] = 16'h0017;
        rom[57][124] = 16'h0008;
        rom[57][125] = 16'h0029;
        rom[57][126] = 16'h000B;
        rom[57][127] = 16'h0023;
        rom[58][0] = 16'hFFFA;
        rom[58][1] = 16'h000E;
        rom[58][2] = 16'hFFE2;
        rom[58][3] = 16'hFFF5;
        rom[58][4] = 16'hFFBA;
        rom[58][5] = 16'h0001;
        rom[58][6] = 16'hFFED;
        rom[58][7] = 16'hFFEF;
        rom[58][8] = 16'hFFD3;
        rom[58][9] = 16'h0000;
        rom[58][10] = 16'hFFBE;
        rom[58][11] = 16'hFFE8;
        rom[58][12] = 16'h0021;
        rom[58][13] = 16'hFFFC;
        rom[58][14] = 16'hFFDF;
        rom[58][15] = 16'hFFE1;
        rom[58][16] = 16'hFFED;
        rom[58][17] = 16'hFFEF;
        rom[58][18] = 16'hFFE5;
        rom[58][19] = 16'hFFE0;
        rom[58][20] = 16'h0011;
        rom[58][21] = 16'hFFD2;
        rom[58][22] = 16'hFFE8;
        rom[58][23] = 16'hFFDA;
        rom[58][24] = 16'hFFDB;
        rom[58][25] = 16'h000A;
        rom[58][26] = 16'hFFF1;
        rom[58][27] = 16'h0007;
        rom[58][28] = 16'hFFDB;
        rom[58][29] = 16'h0007;
        rom[58][30] = 16'hFFF2;
        rom[58][31] = 16'h0003;
        rom[58][32] = 16'hFFF4;
        rom[58][33] = 16'hFFE1;
        rom[58][34] = 16'hFFF0;
        rom[58][35] = 16'h001D;
        rom[58][36] = 16'h000E;
        rom[58][37] = 16'h0011;
        rom[58][38] = 16'hFFD9;
        rom[58][39] = 16'hFFE3;
        rom[58][40] = 16'h0025;
        rom[58][41] = 16'hFFDD;
        rom[58][42] = 16'h0002;
        rom[58][43] = 16'hFFEA;
        rom[58][44] = 16'hFFEF;
        rom[58][45] = 16'h0017;
        rom[58][46] = 16'h0002;
        rom[58][47] = 16'hFFFC;
        rom[58][48] = 16'h001D;
        rom[58][49] = 16'h0017;
        rom[58][50] = 16'hFFEF;
        rom[58][51] = 16'h0015;
        rom[58][52] = 16'h0001;
        rom[58][53] = 16'h001A;
        rom[58][54] = 16'hFFE0;
        rom[58][55] = 16'h001A;
        rom[58][56] = 16'hFFFA;
        rom[58][57] = 16'h0016;
        rom[58][58] = 16'hFFFD;
        rom[58][59] = 16'hFFCF;
        rom[58][60] = 16'hFFD0;
        rom[58][61] = 16'hFFF9;
        rom[58][62] = 16'h0008;
        rom[58][63] = 16'hFFF8;
        rom[58][64] = 16'hFFC6;
        rom[58][65] = 16'h000E;
        rom[58][66] = 16'hFFEA;
        rom[58][67] = 16'h001C;
        rom[58][68] = 16'hFFFF;
        rom[58][69] = 16'h002E;
        rom[58][70] = 16'h0017;
        rom[58][71] = 16'hFFF8;
        rom[58][72] = 16'hFFD2;
        rom[58][73] = 16'h001A;
        rom[58][74] = 16'h0007;
        rom[58][75] = 16'hFFCD;
        rom[58][76] = 16'h001E;
        rom[58][77] = 16'hFFED;
        rom[58][78] = 16'hFFD9;
        rom[58][79] = 16'h0008;
        rom[58][80] = 16'h001D;
        rom[58][81] = 16'hFFEF;
        rom[58][82] = 16'h0017;
        rom[58][83] = 16'hFFE1;
        rom[58][84] = 16'hFFF0;
        rom[58][85] = 16'hFFC7;
        rom[58][86] = 16'hFFD6;
        rom[58][87] = 16'h0010;
        rom[58][88] = 16'hFFEA;
        rom[58][89] = 16'h0021;
        rom[58][90] = 16'h0004;
        rom[58][91] = 16'h0016;
        rom[58][92] = 16'hFFE6;
        rom[58][93] = 16'hFFE6;
        rom[58][94] = 16'h0024;
        rom[58][95] = 16'h0011;
        rom[58][96] = 16'h0001;
        rom[58][97] = 16'h0016;
        rom[58][98] = 16'hFFF0;
        rom[58][99] = 16'hFFF0;
        rom[58][100] = 16'h000C;
        rom[58][101] = 16'hFFD4;
        rom[58][102] = 16'h0018;
        rom[58][103] = 16'h000B;
        rom[58][104] = 16'h0037;
        rom[58][105] = 16'hFFEE;
        rom[58][106] = 16'h000E;
        rom[58][107] = 16'h001D;
        rom[58][108] = 16'hFFC5;
        rom[58][109] = 16'hFFF2;
        rom[58][110] = 16'h001A;
        rom[58][111] = 16'h000E;
        rom[58][112] = 16'h0009;
        rom[58][113] = 16'hFFCD;
        rom[58][114] = 16'h002A;
        rom[58][115] = 16'hFFE5;
        rom[58][116] = 16'hFFFE;
        rom[58][117] = 16'hFFE2;
        rom[58][118] = 16'hFFF1;
        rom[58][119] = 16'hFFF4;
        rom[58][120] = 16'hFFDD;
        rom[58][121] = 16'hFFE3;
        rom[58][122] = 16'hFFF3;
        rom[58][123] = 16'hFFBE;
        rom[58][124] = 16'hFFED;
        rom[58][125] = 16'h0006;
        rom[58][126] = 16'h0016;
        rom[58][127] = 16'hFFFA;
        rom[59][0] = 16'hFFF4;
        rom[59][1] = 16'h000F;
        rom[59][2] = 16'h0004;
        rom[59][3] = 16'hFFFF;
        rom[59][4] = 16'h0022;
        rom[59][5] = 16'h000C;
        rom[59][6] = 16'h002B;
        rom[59][7] = 16'h002D;
        rom[59][8] = 16'h0016;
        rom[59][9] = 16'hFFE6;
        rom[59][10] = 16'hFFEC;
        rom[59][11] = 16'hFFF4;
        rom[59][12] = 16'hFFDD;
        rom[59][13] = 16'h002F;
        rom[59][14] = 16'hFFEC;
        rom[59][15] = 16'h000F;
        rom[59][16] = 16'hFFF4;
        rom[59][17] = 16'h001B;
        rom[59][18] = 16'hFFFA;
        rom[59][19] = 16'hFFC6;
        rom[59][20] = 16'hFFF7;
        rom[59][21] = 16'h0007;
        rom[59][22] = 16'h0015;
        rom[59][23] = 16'h001B;
        rom[59][24] = 16'h0007;
        rom[59][25] = 16'h0005;
        rom[59][26] = 16'hFFF4;
        rom[59][27] = 16'hFFEC;
        rom[59][28] = 16'hFFDC;
        rom[59][29] = 16'hFFD5;
        rom[59][30] = 16'h000E;
        rom[59][31] = 16'h0028;
        rom[59][32] = 16'hFFFE;
        rom[59][33] = 16'h0024;
        rom[59][34] = 16'h0037;
        rom[59][35] = 16'hFFE9;
        rom[59][36] = 16'h002E;
        rom[59][37] = 16'hFFF4;
        rom[59][38] = 16'h000C;
        rom[59][39] = 16'hFFEB;
        rom[59][40] = 16'h0019;
        rom[59][41] = 16'hFFBA;
        rom[59][42] = 16'hFFFF;
        rom[59][43] = 16'hFFF1;
        rom[59][44] = 16'hFFD7;
        rom[59][45] = 16'hFFDF;
        rom[59][46] = 16'h0016;
        rom[59][47] = 16'h0008;
        rom[59][48] = 16'hFFF6;
        rom[59][49] = 16'h0019;
        rom[59][50] = 16'h000D;
        rom[59][51] = 16'h0012;
        rom[59][52] = 16'hFFF0;
        rom[59][53] = 16'hFFEF;
        rom[59][54] = 16'hFFD4;
        rom[59][55] = 16'h0002;
        rom[59][56] = 16'h0003;
        rom[59][57] = 16'h0005;
        rom[59][58] = 16'h000D;
        rom[59][59] = 16'hFFE3;
        rom[59][60] = 16'h000E;
        rom[59][61] = 16'hFFFD;
        rom[59][62] = 16'h0012;
        rom[59][63] = 16'h001B;
        rom[59][64] = 16'h001A;
        rom[59][65] = 16'h0040;
        rom[59][66] = 16'hFFDA;
        rom[59][67] = 16'hFFE0;
        rom[59][68] = 16'h0019;
        rom[59][69] = 16'hFFE5;
        rom[59][70] = 16'h0024;
        rom[59][71] = 16'hFFE2;
        rom[59][72] = 16'hFFF3;
        rom[59][73] = 16'h0002;
        rom[59][74] = 16'hFFFC;
        rom[59][75] = 16'hFFD7;
        rom[59][76] = 16'hFFC1;
        rom[59][77] = 16'hFFC8;
        rom[59][78] = 16'hFFDE;
        rom[59][79] = 16'hFFD0;
        rom[59][80] = 16'hFFF4;
        rom[59][81] = 16'h0004;
        rom[59][82] = 16'h0005;
        rom[59][83] = 16'hFFC6;
        rom[59][84] = 16'h002D;
        rom[59][85] = 16'h0021;
        rom[59][86] = 16'hFFE1;
        rom[59][87] = 16'hFFF4;
        rom[59][88] = 16'h0024;
        rom[59][89] = 16'hFFD7;
        rom[59][90] = 16'hFFF0;
        rom[59][91] = 16'hFFD7;
        rom[59][92] = 16'hFFF3;
        rom[59][93] = 16'hFFCD;
        rom[59][94] = 16'h0012;
        rom[59][95] = 16'h001F;
        rom[59][96] = 16'hFFF6;
        rom[59][97] = 16'hFFE1;
        rom[59][98] = 16'hFFE0;
        rom[59][99] = 16'h0002;
        rom[59][100] = 16'hFFF5;
        rom[59][101] = 16'hFFC8;
        rom[59][102] = 16'hFFEF;
        rom[59][103] = 16'h0033;
        rom[59][104] = 16'h0013;
        rom[59][105] = 16'hFFC3;
        rom[59][106] = 16'hFFEA;
        rom[59][107] = 16'hFFDA;
        rom[59][108] = 16'hFFDC;
        rom[59][109] = 16'h000B;
        rom[59][110] = 16'h001E;
        rom[59][111] = 16'hFFD6;
        rom[59][112] = 16'hFFF2;
        rom[59][113] = 16'hFFE1;
        rom[59][114] = 16'h0021;
        rom[59][115] = 16'h0032;
        rom[59][116] = 16'h001D;
        rom[59][117] = 16'hFFE1;
        rom[59][118] = 16'h0012;
        rom[59][119] = 16'hFFFE;
        rom[59][120] = 16'hFFE0;
        rom[59][121] = 16'hFFF4;
        rom[59][122] = 16'hFFB2;
        rom[59][123] = 16'h0012;
        rom[59][124] = 16'hFFEE;
        rom[59][125] = 16'hFFE8;
        rom[59][126] = 16'hFFEA;
        rom[59][127] = 16'hFFFB;
        rom[60][0] = 16'h0000;
        rom[60][1] = 16'h0026;
        rom[60][2] = 16'h0024;
        rom[60][3] = 16'hFFF0;
        rom[60][4] = 16'h0026;
        rom[60][5] = 16'hFFC5;
        rom[60][6] = 16'h0029;
        rom[60][7] = 16'h0009;
        rom[60][8] = 16'hFFCB;
        rom[60][9] = 16'hFFE1;
        rom[60][10] = 16'hFFEB;
        rom[60][11] = 16'hFFFD;
        rom[60][12] = 16'hFFB4;
        rom[60][13] = 16'hFFFD;
        rom[60][14] = 16'hFFF9;
        rom[60][15] = 16'h0007;
        rom[60][16] = 16'h0002;
        rom[60][17] = 16'h0001;
        rom[60][18] = 16'h0010;
        rom[60][19] = 16'hFFEF;
        rom[60][20] = 16'h0011;
        rom[60][21] = 16'hFFEF;
        rom[60][22] = 16'h0006;
        rom[60][23] = 16'hFFC1;
        rom[60][24] = 16'hFFFA;
        rom[60][25] = 16'hFFB9;
        rom[60][26] = 16'h0005;
        rom[60][27] = 16'hFFF9;
        rom[60][28] = 16'hFFF0;
        rom[60][29] = 16'h0005;
        rom[60][30] = 16'hFFE4;
        rom[60][31] = 16'hFFDA;
        rom[60][32] = 16'h0028;
        rom[60][33] = 16'h0017;
        rom[60][34] = 16'h0024;
        rom[60][35] = 16'hFFEA;
        rom[60][36] = 16'hFFF4;
        rom[60][37] = 16'h0007;
        rom[60][38] = 16'h0004;
        rom[60][39] = 16'hFFFF;
        rom[60][40] = 16'hFFE4;
        rom[60][41] = 16'hFFC9;
        rom[60][42] = 16'hFFA0;
        rom[60][43] = 16'hFFDC;
        rom[60][44] = 16'hFFE9;
        rom[60][45] = 16'h0004;
        rom[60][46] = 16'h0018;
        rom[60][47] = 16'hFFCC;
        rom[60][48] = 16'hFFE3;
        rom[60][49] = 16'hFFD6;
        rom[60][50] = 16'h0024;
        rom[60][51] = 16'hFFDB;
        rom[60][52] = 16'hFFF8;
        rom[60][53] = 16'h0014;
        rom[60][54] = 16'h004F;
        rom[60][55] = 16'hFFB7;
        rom[60][56] = 16'hFFF1;
        rom[60][57] = 16'hFFD0;
        rom[60][58] = 16'h000F;
        rom[60][59] = 16'h000A;
        rom[60][60] = 16'h000C;
        rom[60][61] = 16'hFFD0;
        rom[60][62] = 16'h0004;
        rom[60][63] = 16'h0004;
        rom[60][64] = 16'h003D;
        rom[60][65] = 16'h000C;
        rom[60][66] = 16'h0002;
        rom[60][67] = 16'hFFF5;
        rom[60][68] = 16'h0010;
        rom[60][69] = 16'hFFBA;
        rom[60][70] = 16'hFFF4;
        rom[60][71] = 16'h002C;
        rom[60][72] = 16'hFFFF;
        rom[60][73] = 16'h000C;
        rom[60][74] = 16'hFFF1;
        rom[60][75] = 16'h001E;
        rom[60][76] = 16'hFFDF;
        rom[60][77] = 16'h0011;
        rom[60][78] = 16'h000D;
        rom[60][79] = 16'hFFFD;
        rom[60][80] = 16'h0001;
        rom[60][81] = 16'h003B;
        rom[60][82] = 16'hFFD2;
        rom[60][83] = 16'hFFBF;
        rom[60][84] = 16'h0002;
        rom[60][85] = 16'h0011;
        rom[60][86] = 16'h000C;
        rom[60][87] = 16'h002D;
        rom[60][88] = 16'h0036;
        rom[60][89] = 16'h003E;
        rom[60][90] = 16'hFFEF;
        rom[60][91] = 16'h0004;
        rom[60][92] = 16'h0020;
        rom[60][93] = 16'hFFDF;
        rom[60][94] = 16'h001C;
        rom[60][95] = 16'hFFCF;
        rom[60][96] = 16'hFFF3;
        rom[60][97] = 16'h0012;
        rom[60][98] = 16'hFFBE;
        rom[60][99] = 16'h0019;
        rom[60][100] = 16'hFFC5;
        rom[60][101] = 16'hFFFB;
        rom[60][102] = 16'hFFEA;
        rom[60][103] = 16'hFFF5;
        rom[60][104] = 16'h0005;
        rom[60][105] = 16'hFFE9;
        rom[60][106] = 16'hFFF5;
        rom[60][107] = 16'hFFEB;
        rom[60][108] = 16'h000C;
        rom[60][109] = 16'hFFE2;
        rom[60][110] = 16'hFFFD;
        rom[60][111] = 16'hFFF3;
        rom[60][112] = 16'hFFB5;
        rom[60][113] = 16'h001B;
        rom[60][114] = 16'hFFD2;
        rom[60][115] = 16'hFFF9;
        rom[60][116] = 16'hFFF9;
        rom[60][117] = 16'hFFD2;
        rom[60][118] = 16'hFFFB;
        rom[60][119] = 16'h0004;
        rom[60][120] = 16'hFFF5;
        rom[60][121] = 16'hFFD5;
        rom[60][122] = 16'h001A;
        rom[60][123] = 16'hFFF9;
        rom[60][124] = 16'h0028;
        rom[60][125] = 16'hFFFD;
        rom[60][126] = 16'h001D;
        rom[60][127] = 16'h000C;
        rom[61][0] = 16'hFFFE;
        rom[61][1] = 16'h001E;
        rom[61][2] = 16'hFFDD;
        rom[61][3] = 16'h000E;
        rom[61][4] = 16'hFFE1;
        rom[61][5] = 16'h0017;
        rom[61][6] = 16'hFFDC;
        rom[61][7] = 16'h0006;
        rom[61][8] = 16'h0020;
        rom[61][9] = 16'h0007;
        rom[61][10] = 16'hFFF9;
        rom[61][11] = 16'hFF9F;
        rom[61][12] = 16'h000B;
        rom[61][13] = 16'h0022;
        rom[61][14] = 16'hFFED;
        rom[61][15] = 16'h0004;
        rom[61][16] = 16'hFFDC;
        rom[61][17] = 16'h000D;
        rom[61][18] = 16'hFFF3;
        rom[61][19] = 16'h001B;
        rom[61][20] = 16'hFFEF;
        rom[61][21] = 16'h0004;
        rom[61][22] = 16'hFFFF;
        rom[61][23] = 16'h0020;
        rom[61][24] = 16'hFFEC;
        rom[61][25] = 16'h000D;
        rom[61][26] = 16'hFFE4;
        rom[61][27] = 16'hFFD1;
        rom[61][28] = 16'hFFF9;
        rom[61][29] = 16'h0006;
        rom[61][30] = 16'h0022;
        rom[61][31] = 16'hFFFE;
        rom[61][32] = 16'h000F;
        rom[61][33] = 16'hFFF5;
        rom[61][34] = 16'hFFCE;
        rom[61][35] = 16'hFFD4;
        rom[61][36] = 16'hFFF4;
        rom[61][37] = 16'hFFBC;
        rom[61][38] = 16'h0010;
        rom[61][39] = 16'h0003;
        rom[61][40] = 16'h000D;
        rom[61][41] = 16'hFFF9;
        rom[61][42] = 16'h0001;
        rom[61][43] = 16'hFFE7;
        rom[61][44] = 16'h0008;
        rom[61][45] = 16'hFFD5;
        rom[61][46] = 16'h000C;
        rom[61][47] = 16'hFFE0;
        rom[61][48] = 16'hFFEC;
        rom[61][49] = 16'h0000;
        rom[61][50] = 16'hFFE4;
        rom[61][51] = 16'h0025;
        rom[61][52] = 16'hFFBD;
        rom[61][53] = 16'h0029;
        rom[61][54] = 16'h0029;
        rom[61][55] = 16'hFFFB;
        rom[61][56] = 16'hFFE1;
        rom[61][57] = 16'hFFF4;
        rom[61][58] = 16'hFFF9;
        rom[61][59] = 16'h001B;
        rom[61][60] = 16'h0006;
        rom[61][61] = 16'hFFEE;
        rom[61][62] = 16'h0002;
        rom[61][63] = 16'hFFF0;
        rom[61][64] = 16'h0025;
        rom[61][65] = 16'h000C;
        rom[61][66] = 16'h0014;
        rom[61][67] = 16'h002A;
        rom[61][68] = 16'h002E;
        rom[61][69] = 16'h0021;
        rom[61][70] = 16'hFFE8;
        rom[61][71] = 16'hFFC9;
        rom[61][72] = 16'hFFB1;
        rom[61][73] = 16'h0018;
        rom[61][74] = 16'h001B;
        rom[61][75] = 16'h000F;
        rom[61][76] = 16'hFFB1;
        rom[61][77] = 16'h000C;
        rom[61][78] = 16'h0017;
        rom[61][79] = 16'h0006;
        rom[61][80] = 16'h000E;
        rom[61][81] = 16'hFFFE;
        rom[61][82] = 16'h0011;
        rom[61][83] = 16'h0005;
        rom[61][84] = 16'h000F;
        rom[61][85] = 16'h002E;
        rom[61][86] = 16'h0008;
        rom[61][87] = 16'hFFFC;
        rom[61][88] = 16'h0010;
        rom[61][89] = 16'h001D;
        rom[61][90] = 16'hFFFC;
        rom[61][91] = 16'hFFF5;
        rom[61][92] = 16'hFFE8;
        rom[61][93] = 16'hFFE3;
        rom[61][94] = 16'h000C;
        rom[61][95] = 16'h0004;
        rom[61][96] = 16'h000B;
        rom[61][97] = 16'hFFEE;
        rom[61][98] = 16'hFFE9;
        rom[61][99] = 16'hFFEE;
        rom[61][100] = 16'hFFC7;
        rom[61][101] = 16'hFFE2;
        rom[61][102] = 16'hFFBE;
        rom[61][103] = 16'h0007;
        rom[61][104] = 16'h0028;
        rom[61][105] = 16'hFFFC;
        rom[61][106] = 16'h0009;
        rom[61][107] = 16'hFFC2;
        rom[61][108] = 16'hFFD4;
        rom[61][109] = 16'hFFD5;
        rom[61][110] = 16'h0019;
        rom[61][111] = 16'hFFFD;
        rom[61][112] = 16'h001C;
        rom[61][113] = 16'h0012;
        rom[61][114] = 16'hFFBF;
        rom[61][115] = 16'hFFF9;
        rom[61][116] = 16'h0008;
        rom[61][117] = 16'hFFFE;
        rom[61][118] = 16'h0024;
        rom[61][119] = 16'h0027;
        rom[61][120] = 16'h001A;
        rom[61][121] = 16'h0011;
        rom[61][122] = 16'hFFE6;
        rom[61][123] = 16'h0006;
        rom[61][124] = 16'h0016;
        rom[61][125] = 16'h001F;
        rom[61][126] = 16'hFFC8;
        rom[61][127] = 16'hFFBC;
        rom[62][0] = 16'hFFF5;
        rom[62][1] = 16'hFFCD;
        rom[62][2] = 16'h000B;
        rom[62][3] = 16'h000C;
        rom[62][4] = 16'h0011;
        rom[62][5] = 16'hFFFC;
        rom[62][6] = 16'hFFF9;
        rom[62][7] = 16'hFFC8;
        rom[62][8] = 16'hFFEA;
        rom[62][9] = 16'hFFFE;
        rom[62][10] = 16'hFFE4;
        rom[62][11] = 16'hFFF9;
        rom[62][12] = 16'hFFFD;
        rom[62][13] = 16'hFFD5;
        rom[62][14] = 16'hFFF8;
        rom[62][15] = 16'h0007;
        rom[62][16] = 16'h000F;
        rom[62][17] = 16'hFFF4;
        rom[62][18] = 16'hFFF1;
        rom[62][19] = 16'hFFF2;
        rom[62][20] = 16'h0022;
        rom[62][21] = 16'hFFE6;
        rom[62][22] = 16'h001B;
        rom[62][23] = 16'hFFE6;
        rom[62][24] = 16'h0004;
        rom[62][25] = 16'hFFFE;
        rom[62][26] = 16'hFFFB;
        rom[62][27] = 16'h0034;
        rom[62][28] = 16'h000C;
        rom[62][29] = 16'h0003;
        rom[62][30] = 16'hFFD7;
        rom[62][31] = 16'h0010;
        rom[62][32] = 16'hFFF0;
        rom[62][33] = 16'hFFF4;
        rom[62][34] = 16'h0002;
        rom[62][35] = 16'hFFFC;
        rom[62][36] = 16'hFFCF;
        rom[62][37] = 16'h000A;
        rom[62][38] = 16'h001F;
        rom[62][39] = 16'hFFFA;
        rom[62][40] = 16'hFFE8;
        rom[62][41] = 16'hFFFB;
        rom[62][42] = 16'hFFFC;
        rom[62][43] = 16'h0009;
        rom[62][44] = 16'h000F;
        rom[62][45] = 16'hFFCC;
        rom[62][46] = 16'hFFF2;
        rom[62][47] = 16'h000F;
        rom[62][48] = 16'h000D;
        rom[62][49] = 16'hFFF6;
        rom[62][50] = 16'hFFEF;
        rom[62][51] = 16'h0001;
        rom[62][52] = 16'hFFFB;
        rom[62][53] = 16'hFFE6;
        rom[62][54] = 16'hFFB5;
        rom[62][55] = 16'hFFFB;
        rom[62][56] = 16'hFFE5;
        rom[62][57] = 16'hFFF9;
        rom[62][58] = 16'hFFC8;
        rom[62][59] = 16'h0024;
        rom[62][60] = 16'h0005;
        rom[62][61] = 16'h0011;
        rom[62][62] = 16'hFFFD;
        rom[62][63] = 16'hFFE0;
        rom[62][64] = 16'h0008;
        rom[62][65] = 16'hFFE6;
        rom[62][66] = 16'hFFF3;
        rom[62][67] = 16'hFFF4;
        rom[62][68] = 16'hFFF3;
        rom[62][69] = 16'hFFEC;
        rom[62][70] = 16'h001D;
        rom[62][71] = 16'hFFF1;
        rom[62][72] = 16'hFFF3;
        rom[62][73] = 16'hFFE1;
        rom[62][74] = 16'hFFBA;
        rom[62][75] = 16'hFFF7;
        rom[62][76] = 16'h0003;
        rom[62][77] = 16'hFFEA;
        rom[62][78] = 16'hFFDE;
        rom[62][79] = 16'h0002;
        rom[62][80] = 16'h000D;
        rom[62][81] = 16'hFFC8;
        rom[62][82] = 16'hFFFF;
        rom[62][83] = 16'hFFE5;
        rom[62][84] = 16'h0010;
        rom[62][85] = 16'h001C;
        rom[62][86] = 16'hFFE5;
        rom[62][87] = 16'h0023;
        rom[62][88] = 16'h000A;
        rom[62][89] = 16'hFFE2;
        rom[62][90] = 16'hFFFB;
        rom[62][91] = 16'h0004;
        rom[62][92] = 16'hFFCD;
        rom[62][93] = 16'hFFE8;
        rom[62][94] = 16'hFFEB;
        rom[62][95] = 16'hFFF0;
        rom[62][96] = 16'h0007;
        rom[62][97] = 16'h0014;
        rom[62][98] = 16'hFFEA;
        rom[62][99] = 16'hFFE5;
        rom[62][100] = 16'hFFF4;
        rom[62][101] = 16'hFFFE;
        rom[62][102] = 16'h0011;
        rom[62][103] = 16'h001C;
        rom[62][104] = 16'h001B;
        rom[62][105] = 16'h0000;
        rom[62][106] = 16'h0032;
        rom[62][107] = 16'hFFE0;
        rom[62][108] = 16'hFFE4;
        rom[62][109] = 16'h0041;
        rom[62][110] = 16'h0020;
        rom[62][111] = 16'hFFCE;
        rom[62][112] = 16'h0002;
        rom[62][113] = 16'hFFCB;
        rom[62][114] = 16'h003D;
        rom[62][115] = 16'h0017;
        rom[62][116] = 16'hFFE8;
        rom[62][117] = 16'hFFFC;
        rom[62][118] = 16'hFFF1;
        rom[62][119] = 16'h001D;
        rom[62][120] = 16'hFFF5;
        rom[62][121] = 16'hFFF6;
        rom[62][122] = 16'h0002;
        rom[62][123] = 16'hFFFE;
        rom[62][124] = 16'h0002;
        rom[62][125] = 16'h003A;
        rom[62][126] = 16'h0014;
        rom[62][127] = 16'hFFC7;
        rom[63][0] = 16'hFFD2;
        rom[63][1] = 16'hFFF7;
        rom[63][2] = 16'hFFDE;
        rom[63][3] = 16'hFFFA;
        rom[63][4] = 16'hFFED;
        rom[63][5] = 16'h0032;
        rom[63][6] = 16'h0018;
        rom[63][7] = 16'hFFE6;
        rom[63][8] = 16'h000F;
        rom[63][9] = 16'hFFEE;
        rom[63][10] = 16'h0005;
        rom[63][11] = 16'hFFCF;
        rom[63][12] = 16'hFFF9;
        rom[63][13] = 16'h0004;
        rom[63][14] = 16'h0026;
        rom[63][15] = 16'hFFED;
        rom[63][16] = 16'h001E;
        rom[63][17] = 16'h001B;
        rom[63][18] = 16'hFFE0;
        rom[63][19] = 16'h002D;
        rom[63][20] = 16'hFFFB;
        rom[63][21] = 16'hFFDA;
        rom[63][22] = 16'hFFFE;
        rom[63][23] = 16'hFFF1;
        rom[63][24] = 16'hFFDD;
        rom[63][25] = 16'h000D;
        rom[63][26] = 16'hFFEE;
        rom[63][27] = 16'hFFF3;
        rom[63][28] = 16'hFFEF;
        rom[63][29] = 16'hFFF1;
        rom[63][30] = 16'hFFFC;
        rom[63][31] = 16'h0011;
        rom[63][32] = 16'h001B;
        rom[63][33] = 16'hFFA6;
        rom[63][34] = 16'h000F;
        rom[63][35] = 16'hFFD6;
        rom[63][36] = 16'hFFD3;
        rom[63][37] = 16'hFFE7;
        rom[63][38] = 16'hFFD6;
        rom[63][39] = 16'hFFF7;
        rom[63][40] = 16'hFFF2;
        rom[63][41] = 16'hFFE2;
        rom[63][42] = 16'hFFFE;
        rom[63][43] = 16'hFFC8;
        rom[63][44] = 16'h0019;
        rom[63][45] = 16'hFFF4;
        rom[63][46] = 16'hFFD9;
        rom[63][47] = 16'hFFDE;
        rom[63][48] = 16'hFFFD;
        rom[63][49] = 16'h000A;
        rom[63][50] = 16'h0027;
        rom[63][51] = 16'h0002;
        rom[63][52] = 16'h002F;
        rom[63][53] = 16'h0025;
        rom[63][54] = 16'h0008;
        rom[63][55] = 16'hFFF2;
        rom[63][56] = 16'hFFD9;
        rom[63][57] = 16'h000C;
        rom[63][58] = 16'hFFC3;
        rom[63][59] = 16'hFFF7;
        rom[63][60] = 16'hFFFA;
        rom[63][61] = 16'hFFE7;
        rom[63][62] = 16'hFFF9;
        rom[63][63] = 16'hFFFB;
        rom[63][64] = 16'h0066;
        rom[63][65] = 16'hFFCC;
        rom[63][66] = 16'hFFE5;
        rom[63][67] = 16'h001A;
        rom[63][68] = 16'hFFDA;
        rom[63][69] = 16'h000D;
        rom[63][70] = 16'hFFF7;
        rom[63][71] = 16'h001B;
        rom[63][72] = 16'hFFC3;
        rom[63][73] = 16'hFFD7;
        rom[63][74] = 16'hFFF4;
        rom[63][75] = 16'hFFCB;
        rom[63][76] = 16'hFFC7;
        rom[63][77] = 16'h0022;
        rom[63][78] = 16'h0028;
        rom[63][79] = 16'hFFED;
        rom[63][80] = 16'h0009;
        rom[63][81] = 16'hFFDC;
        rom[63][82] = 16'h000C;
        rom[63][83] = 16'hFFE0;
        rom[63][84] = 16'h0004;
        rom[63][85] = 16'h0029;
        rom[63][86] = 16'hFFFD;
        rom[63][87] = 16'h0002;
        rom[63][88] = 16'h0017;
        rom[63][89] = 16'h000F;
        rom[63][90] = 16'h0006;
        rom[63][91] = 16'h0003;
        rom[63][92] = 16'hFFE2;
        rom[63][93] = 16'hFFE9;
        rom[63][94] = 16'h001D;
        rom[63][95] = 16'hFFD0;
        rom[63][96] = 16'h0009;
        rom[63][97] = 16'h0004;
        rom[63][98] = 16'h0024;
        rom[63][99] = 16'hFFEF;
        rom[63][100] = 16'hFFE4;
        rom[63][101] = 16'hFFCD;
        rom[63][102] = 16'hFFEB;
        rom[63][103] = 16'hFFC9;
        rom[63][104] = 16'hFFFF;
        rom[63][105] = 16'hFFD2;
        rom[63][106] = 16'hFFE7;
        rom[63][107] = 16'h0008;
        rom[63][108] = 16'h001C;
        rom[63][109] = 16'hFFD0;
        rom[63][110] = 16'hFFF7;
        rom[63][111] = 16'hFFF4;
        rom[63][112] = 16'h002E;
        rom[63][113] = 16'hFFF9;
        rom[63][114] = 16'h001C;
        rom[63][115] = 16'hFFE1;
        rom[63][116] = 16'hFFC5;
        rom[63][117] = 16'h0013;
        rom[63][118] = 16'hFFFE;
        rom[63][119] = 16'hFFE4;
        rom[63][120] = 16'hFFDE;
        rom[63][121] = 16'h002B;
        rom[63][122] = 16'hFFE1;
        rom[63][123] = 16'h0018;
        rom[63][124] = 16'hFFF3;
        rom[63][125] = 16'h000A;
        rom[63][126] = 16'h002C;
        rom[63][127] = 16'h0025;
        rom[64][0] = 16'hFFF6;
        rom[64][1] = 16'h001A;
        rom[64][2] = 16'hFFDB;
        rom[64][3] = 16'hFFF8;
        rom[64][4] = 16'hFFF4;
        rom[64][5] = 16'h0000;
        rom[64][6] = 16'h0006;
        rom[64][7] = 16'h0038;
        rom[64][8] = 16'h0014;
        rom[64][9] = 16'hFFCF;
        rom[64][10] = 16'hFFD9;
        rom[64][11] = 16'hFFE6;
        rom[64][12] = 16'h0010;
        rom[64][13] = 16'h004D;
        rom[64][14] = 16'hFFF1;
        rom[64][15] = 16'h0007;
        rom[64][16] = 16'h0002;
        rom[64][17] = 16'h0031;
        rom[64][18] = 16'hFFE3;
        rom[64][19] = 16'h0018;
        rom[64][20] = 16'hFFCD;
        rom[64][21] = 16'h0025;
        rom[64][22] = 16'h0011;
        rom[64][23] = 16'hFFB5;
        rom[64][24] = 16'hFFF5;
        rom[64][25] = 16'h0026;
        rom[64][26] = 16'h000A;
        rom[64][27] = 16'hFFD4;
        rom[64][28] = 16'h0014;
        rom[64][29] = 16'h0031;
        rom[64][30] = 16'h0008;
        rom[64][31] = 16'h0016;
        rom[64][32] = 16'h001C;
        rom[64][33] = 16'h001C;
        rom[64][34] = 16'h0018;
        rom[64][35] = 16'hFFF3;
        rom[64][36] = 16'h0005;
        rom[64][37] = 16'hFFE9;
        rom[64][38] = 16'hFFD0;
        rom[64][39] = 16'hFFF9;
        rom[64][40] = 16'h0005;
        rom[64][41] = 16'hFFF9;
        rom[64][42] = 16'hFFF8;
        rom[64][43] = 16'h001F;
        rom[64][44] = 16'hFFE5;
        rom[64][45] = 16'hFFDA;
        rom[64][46] = 16'hFFE4;
        rom[64][47] = 16'h0011;
        rom[64][48] = 16'hFFFF;
        rom[64][49] = 16'h0028;
        rom[64][50] = 16'hFFD1;
        rom[64][51] = 16'hFFF5;
        rom[64][52] = 16'h001B;
        rom[64][53] = 16'h0009;
        rom[64][54] = 16'h0027;
        rom[64][55] = 16'h0001;
        rom[64][56] = 16'hFFF9;
        rom[64][57] = 16'h0007;
        rom[64][58] = 16'hFFF5;
        rom[64][59] = 16'hFFC6;
        rom[64][60] = 16'hFFF3;
        rom[64][61] = 16'h000D;
        rom[64][62] = 16'h000C;
        rom[64][63] = 16'hFFF5;
        rom[64][64] = 16'h000B;
        rom[64][65] = 16'h002E;
        rom[64][66] = 16'h000C;
        rom[64][67] = 16'h0028;
        rom[64][68] = 16'h0043;
        rom[64][69] = 16'h0025;
        rom[64][70] = 16'hFFF9;
        rom[64][71] = 16'h0003;
        rom[64][72] = 16'hFFFB;
        rom[64][73] = 16'hFFF0;
        rom[64][74] = 16'h0015;
        rom[64][75] = 16'hFFF2;
        rom[64][76] = 16'hFFD8;
        rom[64][77] = 16'hFFB9;
        rom[64][78] = 16'h000D;
        rom[64][79] = 16'h0003;
        rom[64][80] = 16'h0011;
        rom[64][81] = 16'hFFF9;
        rom[64][82] = 16'h001B;
        rom[64][83] = 16'h0012;
        rom[64][84] = 16'h002E;
        rom[64][85] = 16'hFFD2;
        rom[64][86] = 16'hFFEF;
        rom[64][87] = 16'h0007;
        rom[64][88] = 16'hFFED;
        rom[64][89] = 16'h000F;
        rom[64][90] = 16'hFFFF;
        rom[64][91] = 16'h0012;
        rom[64][92] = 16'h0005;
        rom[64][93] = 16'h0001;
        rom[64][94] = 16'h001E;
        rom[64][95] = 16'h0012;
        rom[64][96] = 16'h0030;
        rom[64][97] = 16'h0007;
        rom[64][98] = 16'hFFED;
        rom[64][99] = 16'hFFEA;
        rom[64][100] = 16'hFFF2;
        rom[64][101] = 16'hFFC8;
        rom[64][102] = 16'h0001;
        rom[64][103] = 16'hFFDE;
        rom[64][104] = 16'hFFFB;
        rom[64][105] = 16'hFFF8;
        rom[64][106] = 16'hFFE8;
        rom[64][107] = 16'hFFDC;
        rom[64][108] = 16'h0030;
        rom[64][109] = 16'hFFF2;
        rom[64][110] = 16'hFFF4;
        rom[64][111] = 16'hFFCC;
        rom[64][112] = 16'hFFF9;
        rom[64][113] = 16'h0024;
        rom[64][114] = 16'hFFFF;
        rom[64][115] = 16'h000C;
        rom[64][116] = 16'h002A;
        rom[64][117] = 16'h000A;
        rom[64][118] = 16'hFFC6;
        rom[64][119] = 16'hFFE7;
        rom[64][120] = 16'hFFE5;
        rom[64][121] = 16'hFFD3;
        rom[64][122] = 16'hFFCC;
        rom[64][123] = 16'hFFD9;
        rom[64][124] = 16'h0007;
        rom[64][125] = 16'hFFCD;
        rom[64][126] = 16'hFFDE;
        rom[64][127] = 16'hFFEF;
        rom[65][0] = 16'hFFCB;
        rom[65][1] = 16'h0025;
        rom[65][2] = 16'hFFD7;
        rom[65][3] = 16'hFFFE;
        rom[65][4] = 16'hFFFD;
        rom[65][5] = 16'h0022;
        rom[65][6] = 16'h0002;
        rom[65][7] = 16'h002A;
        rom[65][8] = 16'hFFF8;
        rom[65][9] = 16'h000A;
        rom[65][10] = 16'h000C;
        rom[65][11] = 16'h001E;
        rom[65][12] = 16'hFFE9;
        rom[65][13] = 16'hFFE2;
        rom[65][14] = 16'hFFDC;
        rom[65][15] = 16'h000B;
        rom[65][16] = 16'h001F;
        rom[65][17] = 16'h0009;
        rom[65][18] = 16'h002E;
        rom[65][19] = 16'h0008;
        rom[65][20] = 16'hFFBC;
        rom[65][21] = 16'h002E;
        rom[65][22] = 16'hFFCE;
        rom[65][23] = 16'hFFF7;
        rom[65][24] = 16'hFFEF;
        rom[65][25] = 16'hFFEF;
        rom[65][26] = 16'h001B;
        rom[65][27] = 16'hFFEF;
        rom[65][28] = 16'hFFEA;
        rom[65][29] = 16'h000F;
        rom[65][30] = 16'h0024;
        rom[65][31] = 16'h0005;
        rom[65][32] = 16'hFFF2;
        rom[65][33] = 16'hFFFD;
        rom[65][34] = 16'h0016;
        rom[65][35] = 16'hFFBA;
        rom[65][36] = 16'h0017;
        rom[65][37] = 16'hFFF1;
        rom[65][38] = 16'hFFD1;
        rom[65][39] = 16'hFFDC;
        rom[65][40] = 16'hFFF9;
        rom[65][41] = 16'hFFF5;
        rom[65][42] = 16'h001F;
        rom[65][43] = 16'h000F;
        rom[65][44] = 16'h0002;
        rom[65][45] = 16'h000E;
        rom[65][46] = 16'hFFF8;
        rom[65][47] = 16'h0002;
        rom[65][48] = 16'hFFBA;
        rom[65][49] = 16'hFFE7;
        rom[65][50] = 16'hFFF4;
        rom[65][51] = 16'hFFE1;
        rom[65][52] = 16'h000D;
        rom[65][53] = 16'h0002;
        rom[65][54] = 16'h0007;
        rom[65][55] = 16'hFFFE;
        rom[65][56] = 16'h0007;
        rom[65][57] = 16'hFFDD;
        rom[65][58] = 16'hFFDF;
        rom[65][59] = 16'h0022;
        rom[65][60] = 16'h0010;
        rom[65][61] = 16'h000A;
        rom[65][62] = 16'hFFF1;
        rom[65][63] = 16'hFFD3;
        rom[65][64] = 16'hFFCD;
        rom[65][65] = 16'h0015;
        rom[65][66] = 16'h000B;
        rom[65][67] = 16'h0032;
        rom[65][68] = 16'h0007;
        rom[65][69] = 16'h0047;
        rom[65][70] = 16'h0022;
        rom[65][71] = 16'hFFFD;
        rom[65][72] = 16'hFFF1;
        rom[65][73] = 16'h0024;
        rom[65][74] = 16'hFFEF;
        rom[65][75] = 16'h0002;
        rom[65][76] = 16'hFFF9;
        rom[65][77] = 16'h0019;
        rom[65][78] = 16'h0045;
        rom[65][79] = 16'h0010;
        rom[65][80] = 16'h004A;
        rom[65][81] = 16'h001B;
        rom[65][82] = 16'h0011;
        rom[65][83] = 16'h0015;
        rom[65][84] = 16'h0004;
        rom[65][85] = 16'hFFE1;
        rom[65][86] = 16'hFFF6;
        rom[65][87] = 16'h0002;
        rom[65][88] = 16'hFFD8;
        rom[65][89] = 16'hFFD9;
        rom[65][90] = 16'hFFF5;
        rom[65][91] = 16'h002E;
        rom[65][92] = 16'hFFF6;
        rom[65][93] = 16'h000C;
        rom[65][94] = 16'hFFF9;
        rom[65][95] = 16'hFFE8;
        rom[65][96] = 16'h001B;
        rom[65][97] = 16'hFFDC;
        rom[65][98] = 16'hFFFF;
        rom[65][99] = 16'h000F;
        rom[65][100] = 16'h0019;
        rom[65][101] = 16'hFFDF;
        rom[65][102] = 16'hFFCF;
        rom[65][103] = 16'hFFF9;
        rom[65][104] = 16'h0012;
        rom[65][105] = 16'hFFDE;
        rom[65][106] = 16'h0011;
        rom[65][107] = 16'h004B;
        rom[65][108] = 16'hFFEA;
        rom[65][109] = 16'hFFD3;
        rom[65][110] = 16'hFFE3;
        rom[65][111] = 16'hFFFE;
        rom[65][112] = 16'hFFCC;
        rom[65][113] = 16'hFFC5;
        rom[65][114] = 16'hFFCB;
        rom[65][115] = 16'hFFF1;
        rom[65][116] = 16'h0001;
        rom[65][117] = 16'hFFEA;
        rom[65][118] = 16'hFFD2;
        rom[65][119] = 16'hFFD0;
        rom[65][120] = 16'hFFF3;
        rom[65][121] = 16'hFFCD;
        rom[65][122] = 16'h0022;
        rom[65][123] = 16'hFFEC;
        rom[65][124] = 16'h0012;
        rom[65][125] = 16'h001C;
        rom[65][126] = 16'h0011;
        rom[65][127] = 16'h0003;
        rom[66][0] = 16'h0015;
        rom[66][1] = 16'hFFA3;
        rom[66][2] = 16'h0036;
        rom[66][3] = 16'hFFFE;
        rom[66][4] = 16'h0002;
        rom[66][5] = 16'hFFEB;
        rom[66][6] = 16'h0007;
        rom[66][7] = 16'hFFEE;
        rom[66][8] = 16'hFFE2;
        rom[66][9] = 16'h0002;
        rom[66][10] = 16'h002E;
        rom[66][11] = 16'h0002;
        rom[66][12] = 16'hFFC8;
        rom[66][13] = 16'h001E;
        rom[66][14] = 16'h0006;
        rom[66][15] = 16'h0004;
        rom[66][16] = 16'h002D;
        rom[66][17] = 16'h0010;
        rom[66][18] = 16'h0010;
        rom[66][19] = 16'h000E;
        rom[66][20] = 16'hFFF2;
        rom[66][21] = 16'hFFEB;
        rom[66][22] = 16'h0013;
        rom[66][23] = 16'hFFFA;
        rom[66][24] = 16'hFFDE;
        rom[66][25] = 16'h000A;
        rom[66][26] = 16'h000D;
        rom[66][27] = 16'h0013;
        rom[66][28] = 16'h0024;
        rom[66][29] = 16'hFFF9;
        rom[66][30] = 16'hFFEF;
        rom[66][31] = 16'hFFB2;
        rom[66][32] = 16'h0023;
        rom[66][33] = 16'hFFF7;
        rom[66][34] = 16'hFFFC;
        rom[66][35] = 16'hFFF5;
        rom[66][36] = 16'hFFAE;
        rom[66][37] = 16'hFFE1;
        rom[66][38] = 16'h0016;
        rom[66][39] = 16'hFFE4;
        rom[66][40] = 16'hFFE1;
        rom[66][41] = 16'hFFDF;
        rom[66][42] = 16'h0012;
        rom[66][43] = 16'hFFD7;
        rom[66][44] = 16'hFFEA;
        rom[66][45] = 16'h0013;
        rom[66][46] = 16'hFFDB;
        rom[66][47] = 16'hFFD6;
        rom[66][48] = 16'hFFA8;
        rom[66][49] = 16'h001B;
        rom[66][50] = 16'h000A;
        rom[66][51] = 16'h0029;
        rom[66][52] = 16'h0000;
        rom[66][53] = 16'hFFDA;
        rom[66][54] = 16'hFFD7;
        rom[66][55] = 16'hFFE8;
        rom[66][56] = 16'hFFDC;
        rom[66][57] = 16'h0007;
        rom[66][58] = 16'hFFCC;
        rom[66][59] = 16'h001B;
        rom[66][60] = 16'h001B;
        rom[66][61] = 16'hFFD7;
        rom[66][62] = 16'h001B;
        rom[66][63] = 16'hFFBF;
        rom[66][64] = 16'h0002;
        rom[66][65] = 16'hFFE1;
        rom[66][66] = 16'h000A;
        rom[66][67] = 16'hFFF9;
        rom[66][68] = 16'h0023;
        rom[66][69] = 16'hFFE7;
        rom[66][70] = 16'h0013;
        rom[66][71] = 16'h0011;
        rom[66][72] = 16'hFFCF;
        rom[66][73] = 16'h0001;
        rom[66][74] = 16'hFFD2;
        rom[66][75] = 16'hFFD5;
        rom[66][76] = 16'hFFE1;
        rom[66][77] = 16'hFFFD;
        rom[66][78] = 16'hFFF4;
        rom[66][79] = 16'hFFB5;
        rom[66][80] = 16'hFFE1;
        rom[66][81] = 16'hFFB8;
        rom[66][82] = 16'hFFF1;
        rom[66][83] = 16'hFFE5;
        rom[66][84] = 16'hFFFB;
        rom[66][85] = 16'h0016;
        rom[66][86] = 16'h000F;
        rom[66][87] = 16'h0009;
        rom[66][88] = 16'h001C;
        rom[66][89] = 16'hFFF0;
        rom[66][90] = 16'h0004;
        rom[66][91] = 16'h0034;
        rom[66][92] = 16'h0026;
        rom[66][93] = 16'hFFE5;
        rom[66][94] = 16'h0000;
        rom[66][95] = 16'hFFFF;
        rom[66][96] = 16'hFFDF;
        rom[66][97] = 16'hFFFF;
        rom[66][98] = 16'h000A;
        rom[66][99] = 16'hFFE2;
        rom[66][100] = 16'h0048;
        rom[66][101] = 16'hFFBE;
        rom[66][102] = 16'hFFF3;
        rom[66][103] = 16'hFFC1;
        rom[66][104] = 16'h0013;
        rom[66][105] = 16'hFFD8;
        rom[66][106] = 16'hFFF5;
        rom[66][107] = 16'h0011;
        rom[66][108] = 16'h0033;
        rom[66][109] = 16'h0000;
        rom[66][110] = 16'h0010;
        rom[66][111] = 16'hFFEF;
        rom[66][112] = 16'hFFEA;
        rom[66][113] = 16'h0041;
        rom[66][114] = 16'h000A;
        rom[66][115] = 16'hFFE1;
        rom[66][116] = 16'hFFFE;
        rom[66][117] = 16'h0002;
        rom[66][118] = 16'hFFE1;
        rom[66][119] = 16'hFFFF;
        rom[66][120] = 16'h0012;
        rom[66][121] = 16'h0021;
        rom[66][122] = 16'h0016;
        rom[66][123] = 16'h0038;
        rom[66][124] = 16'h000C;
        rom[66][125] = 16'hFFFC;
        rom[66][126] = 16'h0029;
        rom[66][127] = 16'h0010;
        rom[67][0] = 16'hFFE3;
        rom[67][1] = 16'h0032;
        rom[67][2] = 16'h0009;
        rom[67][3] = 16'h0013;
        rom[67][4] = 16'hFFF5;
        rom[67][5] = 16'h0029;
        rom[67][6] = 16'hFFE7;
        rom[67][7] = 16'hFFF8;
        rom[67][8] = 16'h0002;
        rom[67][9] = 16'hFFF4;
        rom[67][10] = 16'hFFF9;
        rom[67][11] = 16'hFFFD;
        rom[67][12] = 16'h002F;
        rom[67][13] = 16'h0009;
        rom[67][14] = 16'hFFCA;
        rom[67][15] = 16'h0024;
        rom[67][16] = 16'h0002;
        rom[67][17] = 16'h0013;
        rom[67][18] = 16'hFFCD;
        rom[67][19] = 16'h001A;
        rom[67][20] = 16'hFFF2;
        rom[67][21] = 16'h0027;
        rom[67][22] = 16'hFFE8;
        rom[67][23] = 16'hFFF0;
        rom[67][24] = 16'h0003;
        rom[67][25] = 16'h0014;
        rom[67][26] = 16'h0012;
        rom[67][27] = 16'h002D;
        rom[67][28] = 16'h0015;
        rom[67][29] = 16'hFFF9;
        rom[67][30] = 16'h0033;
        rom[67][31] = 16'h0002;
        rom[67][32] = 16'h0006;
        rom[67][33] = 16'hFFFA;
        rom[67][34] = 16'hFFF1;
        rom[67][35] = 16'h0022;
        rom[67][36] = 16'hFFD7;
        rom[67][37] = 16'h002E;
        rom[67][38] = 16'hFFD6;
        rom[67][39] = 16'hFFE0;
        rom[67][40] = 16'h0015;
        rom[67][41] = 16'h0002;
        rom[67][42] = 16'h0010;
        rom[67][43] = 16'hFFEA;
        rom[67][44] = 16'hFFE0;
        rom[67][45] = 16'h001A;
        rom[67][46] = 16'hFFC0;
        rom[67][47] = 16'h0022;
        rom[67][48] = 16'h0007;
        rom[67][49] = 16'hFFF6;
        rom[67][50] = 16'hFFFE;
        rom[67][51] = 16'hFFCD;
        rom[67][52] = 16'hFFF5;
        rom[67][53] = 16'hFFFA;
        rom[67][54] = 16'hFFF5;
        rom[67][55] = 16'h0005;
        rom[67][56] = 16'hFFE3;
        rom[67][57] = 16'hFFDA;
        rom[67][58] = 16'hFFEC;
        rom[67][59] = 16'h0035;
        rom[67][60] = 16'hFFFE;
        rom[67][61] = 16'h0007;
        rom[67][62] = 16'h000C;
        rom[67][63] = 16'h000C;
        rom[67][64] = 16'h0003;
        rom[67][65] = 16'hFFE9;
        rom[67][66] = 16'hFFF7;
        rom[67][67] = 16'h0009;
        rom[67][68] = 16'hFFB9;
        rom[67][69] = 16'h0008;
        rom[67][70] = 16'h0025;
        rom[67][71] = 16'hFFFB;
        rom[67][72] = 16'h000E;
        rom[67][73] = 16'h001C;
        rom[67][74] = 16'hFFD0;
        rom[67][75] = 16'h0011;
        rom[67][76] = 16'hFFE0;
        rom[67][77] = 16'hFFEA;
        rom[67][78] = 16'hFFFE;
        rom[67][79] = 16'hFFF6;
        rom[67][80] = 16'hFFFB;
        rom[67][81] = 16'hFFFE;
        rom[67][82] = 16'h0036;
        rom[67][83] = 16'h0002;
        rom[67][84] = 16'hFFD9;
        rom[67][85] = 16'h0015;
        rom[67][86] = 16'hFFE3;
        rom[67][87] = 16'hFFE9;
        rom[67][88] = 16'hFFE9;
        rom[67][89] = 16'h0015;
        rom[67][90] = 16'h0018;
        rom[67][91] = 16'hFFA8;
        rom[67][92] = 16'h0005;
        rom[67][93] = 16'h0013;
        rom[67][94] = 16'hFFF6;
        rom[67][95] = 16'hFFFB;
        rom[67][96] = 16'hFFDC;
        rom[67][97] = 16'hFFE2;
        rom[67][98] = 16'h0014;
        rom[67][99] = 16'hFFF2;
        rom[67][100] = 16'hFFFF;
        rom[67][101] = 16'h0001;
        rom[67][102] = 16'hFFE4;
        rom[67][103] = 16'hFFD0;
        rom[67][104] = 16'h0007;
        rom[67][105] = 16'h0016;
        rom[67][106] = 16'h0028;
        rom[67][107] = 16'h0007;
        rom[67][108] = 16'hFFF2;
        rom[67][109] = 16'h0023;
        rom[67][110] = 16'h0038;
        rom[67][111] = 16'h0008;
        rom[67][112] = 16'h001D;
        rom[67][113] = 16'hFFEB;
        rom[67][114] = 16'h000D;
        rom[67][115] = 16'hFFF8;
        rom[67][116] = 16'hFFFA;
        rom[67][117] = 16'hFFEF;
        rom[67][118] = 16'h0013;
        rom[67][119] = 16'h000B;
        rom[67][120] = 16'h0007;
        rom[67][121] = 16'hFFFA;
        rom[67][122] = 16'h0000;
        rom[67][123] = 16'hFFE5;
        rom[67][124] = 16'hFFEC;
        rom[67][125] = 16'hFFDF;
        rom[67][126] = 16'h0028;
        rom[67][127] = 16'hFFF8;
        rom[68][0] = 16'h001B;
        rom[68][1] = 16'hFFF9;
        rom[68][2] = 16'h0010;
        rom[68][3] = 16'h0009;
        rom[68][4] = 16'hFFC9;
        rom[68][5] = 16'hFFF0;
        rom[68][6] = 16'h0017;
        rom[68][7] = 16'h0007;
        rom[68][8] = 16'hFFFC;
        rom[68][9] = 16'h0019;
        rom[68][10] = 16'hFFD6;
        rom[68][11] = 16'h0009;
        rom[68][12] = 16'hFFE6;
        rom[68][13] = 16'hFFF3;
        rom[68][14] = 16'hFFF1;
        rom[68][15] = 16'hFFF4;
        rom[68][16] = 16'hFFE2;
        rom[68][17] = 16'h0024;
        rom[68][18] = 16'h0011;
        rom[68][19] = 16'hFFCD;
        rom[68][20] = 16'hFFE2;
        rom[68][21] = 16'hFFF1;
        rom[68][22] = 16'h002D;
        rom[68][23] = 16'hFFD7;
        rom[68][24] = 16'h000B;
        rom[68][25] = 16'hFFF4;
        rom[68][26] = 16'hFFE1;
        rom[68][27] = 16'h0005;
        rom[68][28] = 16'h0016;
        rom[68][29] = 16'h001E;
        rom[68][30] = 16'hFFF2;
        rom[68][31] = 16'h0002;
        rom[68][32] = 16'h0016;
        rom[68][33] = 16'h001D;
        rom[68][34] = 16'hFFF9;
        rom[68][35] = 16'h0018;
        rom[68][36] = 16'hFFF6;
        rom[68][37] = 16'hFFEF;
        rom[68][38] = 16'hFFF1;
        rom[68][39] = 16'h0014;
        rom[68][40] = 16'h0006;
        rom[68][41] = 16'hFFF4;
        rom[68][42] = 16'hFFE7;
        rom[68][43] = 16'hFFFE;
        rom[68][44] = 16'h001E;
        rom[68][45] = 16'h0013;
        rom[68][46] = 16'hFFE3;
        rom[68][47] = 16'hFFDC;
        rom[68][48] = 16'hFFF5;
        rom[68][49] = 16'hFFF2;
        rom[68][50] = 16'h000B;
        rom[68][51] = 16'h000E;
        rom[68][52] = 16'h004A;
        rom[68][53] = 16'h0013;
        rom[68][54] = 16'h000D;
        rom[68][55] = 16'h0002;
        rom[68][56] = 16'hFFF5;
        rom[68][57] = 16'hFFEA;
        rom[68][58] = 16'h0000;
        rom[68][59] = 16'hFFD7;
        rom[68][60] = 16'h0001;
        rom[68][61] = 16'h001D;
        rom[68][62] = 16'h0000;
        rom[68][63] = 16'h0001;
        rom[68][64] = 16'h0025;
        rom[68][65] = 16'hFFF8;
        rom[68][66] = 16'hFFE2;
        rom[68][67] = 16'hFFB2;
        rom[68][68] = 16'hFFF0;
        rom[68][69] = 16'hFFEA;
        rom[68][70] = 16'h0006;
        rom[68][71] = 16'h0031;
        rom[68][72] = 16'hFFDC;
        rom[68][73] = 16'h0009;
        rom[68][74] = 16'h0002;
        rom[68][75] = 16'h001B;
        rom[68][76] = 16'hFFFE;
        rom[68][77] = 16'hFFCB;
        rom[68][78] = 16'hFFFB;
        rom[68][79] = 16'hFFE9;
        rom[68][80] = 16'h000C;
        rom[68][81] = 16'h0011;
        rom[68][82] = 16'hFFE6;
        rom[68][83] = 16'h0004;
        rom[68][84] = 16'h002B;
        rom[68][85] = 16'hFFC2;
        rom[68][86] = 16'hFFFA;
        rom[68][87] = 16'hFFC3;
        rom[68][88] = 16'hFFF5;
        rom[68][89] = 16'hFFD7;
        rom[68][90] = 16'hFFEA;
        rom[68][91] = 16'hFFD7;
        rom[68][92] = 16'h0014;
        rom[68][93] = 16'h0003;
        rom[68][94] = 16'hFFC7;
        rom[68][95] = 16'h001F;
        rom[68][96] = 16'hFFFA;
        rom[68][97] = 16'hFFF4;
        rom[68][98] = 16'hFFEA;
        rom[68][99] = 16'hFFEE;
        rom[68][100] = 16'h0014;
        rom[68][101] = 16'h001F;
        rom[68][102] = 16'h0021;
        rom[68][103] = 16'h001A;
        rom[68][104] = 16'hFFF3;
        rom[68][105] = 16'h001B;
        rom[68][106] = 16'h001A;
        rom[68][107] = 16'hFFED;
        rom[68][108] = 16'h000C;
        rom[68][109] = 16'h001E;
        rom[68][110] = 16'hFFC6;
        rom[68][111] = 16'hFFD8;
        rom[68][112] = 16'hFFDF;
        rom[68][113] = 16'h000F;
        rom[68][114] = 16'hFFFA;
        rom[68][115] = 16'hFFEF;
        rom[68][116] = 16'hFFFD;
        rom[68][117] = 16'hFFE8;
        rom[68][118] = 16'hFFCF;
        rom[68][119] = 16'h0007;
        rom[68][120] = 16'h0029;
        rom[68][121] = 16'hFFC9;
        rom[68][122] = 16'h000E;
        rom[68][123] = 16'h0000;
        rom[68][124] = 16'hFFF9;
        rom[68][125] = 16'hFFDA;
        rom[68][126] = 16'hFFF3;
        rom[68][127] = 16'h0038;
        rom[69][0] = 16'hFFFB;
        rom[69][1] = 16'hFFF4;
        rom[69][2] = 16'h001A;
        rom[69][3] = 16'hFFEB;
        rom[69][4] = 16'hFFF6;
        rom[69][5] = 16'h0000;
        rom[69][6] = 16'h0007;
        rom[69][7] = 16'hFFEF;
        rom[69][8] = 16'h0030;
        rom[69][9] = 16'hFFD2;
        rom[69][10] = 16'hFFEE;
        rom[69][11] = 16'hFFEC;
        rom[69][12] = 16'hFFE5;
        rom[69][13] = 16'h0025;
        rom[69][14] = 16'hFFE1;
        rom[69][15] = 16'hFFF4;
        rom[69][16] = 16'hFFCA;
        rom[69][17] = 16'hFFFF;
        rom[69][18] = 16'h0016;
        rom[69][19] = 16'h001B;
        rom[69][20] = 16'h0028;
        rom[69][21] = 16'hFFF1;
        rom[69][22] = 16'h0005;
        rom[69][23] = 16'hFFD8;
        rom[69][24] = 16'hFFEE;
        rom[69][25] = 16'h0010;
        rom[69][26] = 16'h000C;
        rom[69][27] = 16'h0000;
        rom[69][28] = 16'h001F;
        rom[69][29] = 16'h000A;
        rom[69][30] = 16'hFFDC;
        rom[69][31] = 16'hFFFB;
        rom[69][32] = 16'h0025;
        rom[69][33] = 16'h0001;
        rom[69][34] = 16'h0011;
        rom[69][35] = 16'hFFFD;
        rom[69][36] = 16'hFFB9;
        rom[69][37] = 16'hFFDB;
        rom[69][38] = 16'hFFDC;
        rom[69][39] = 16'h0005;
        rom[69][40] = 16'h0009;
        rom[69][41] = 16'hFFE7;
        rom[69][42] = 16'hFFFC;
        rom[69][43] = 16'h003B;
        rom[69][44] = 16'hFFE1;
        rom[69][45] = 16'h0001;
        rom[69][46] = 16'hFFBE;
        rom[69][47] = 16'h001F;
        rom[69][48] = 16'hFFD2;
        rom[69][49] = 16'hFFD7;
        rom[69][50] = 16'hFFDB;
        rom[69][51] = 16'hFFD7;
        rom[69][52] = 16'hFFFE;
        rom[69][53] = 16'hFFF4;
        rom[69][54] = 16'hFFF7;
        rom[69][55] = 16'h0011;
        rom[69][56] = 16'h0006;
        rom[69][57] = 16'hFFF4;
        rom[69][58] = 16'hFFE7;
        rom[69][59] = 16'h000A;
        rom[69][60] = 16'hFFB0;
        rom[69][61] = 16'h0005;
        rom[69][62] = 16'hFFFC;
        rom[69][63] = 16'hFFEE;
        rom[69][64] = 16'h0012;
        rom[69][65] = 16'hFFD1;
        rom[69][66] = 16'hFFF6;
        rom[69][67] = 16'h0018;
        rom[69][68] = 16'h000D;
        rom[69][69] = 16'h0035;
        rom[69][70] = 16'h0007;
        rom[69][71] = 16'h000A;
        rom[69][72] = 16'hFFF3;
        rom[69][73] = 16'hFFDB;
        rom[69][74] = 16'h0005;
        rom[69][75] = 16'hFFF6;
        rom[69][76] = 16'h000C;
        rom[69][77] = 16'hFFED;
        rom[69][78] = 16'hFFED;
        rom[69][79] = 16'hFFDB;
        rom[69][80] = 16'h0023;
        rom[69][81] = 16'hFFC3;
        rom[69][82] = 16'hFFEA;
        rom[69][83] = 16'h0025;
        rom[69][84] = 16'hFFE3;
        rom[69][85] = 16'hFFE4;
        rom[69][86] = 16'hFFE8;
        rom[69][87] = 16'hFFE3;
        rom[69][88] = 16'h0003;
        rom[69][89] = 16'hFFF6;
        rom[69][90] = 16'h0001;
        rom[69][91] = 16'h000A;
        rom[69][92] = 16'hFFF8;
        rom[69][93] = 16'hFFFA;
        rom[69][94] = 16'hFFF1;
        rom[69][95] = 16'hFFDD;
        rom[69][96] = 16'hFFFD;
        rom[69][97] = 16'hFFF7;
        rom[69][98] = 16'h0013;
        rom[69][99] = 16'hFFD7;
        rom[69][100] = 16'h000C;
        rom[69][101] = 16'h0007;
        rom[69][102] = 16'hFFEB;
        rom[69][103] = 16'hFFEA;
        rom[69][104] = 16'hFFD7;
        rom[69][105] = 16'hFFCD;
        rom[69][106] = 16'hFFE5;
        rom[69][107] = 16'hFFF2;
        rom[69][108] = 16'h000E;
        rom[69][109] = 16'hFFC7;
        rom[69][110] = 16'hFFFE;
        rom[69][111] = 16'h000D;
        rom[69][112] = 16'h001C;
        rom[69][113] = 16'h001A;
        rom[69][114] = 16'hFFE9;
        rom[69][115] = 16'hFFFA;
        rom[69][116] = 16'hFFD1;
        rom[69][117] = 16'hFFE5;
        rom[69][118] = 16'h0016;
        rom[69][119] = 16'hFFAD;
        rom[69][120] = 16'hFFD5;
        rom[69][121] = 16'h000B;
        rom[69][122] = 16'hFFC5;
        rom[69][123] = 16'h0009;
        rom[69][124] = 16'hFFF3;
        rom[69][125] = 16'hFFED;
        rom[69][126] = 16'hFFF7;
        rom[69][127] = 16'h000B;
        rom[70][0] = 16'h0034;
        rom[70][1] = 16'hFFDB;
        rom[70][2] = 16'h000C;
        rom[70][3] = 16'hFFD7;
        rom[70][4] = 16'hFFB5;
        rom[70][5] = 16'hFFD3;
        rom[70][6] = 16'hFFD0;
        rom[70][7] = 16'h000E;
        rom[70][8] = 16'hFFC2;
        rom[70][9] = 16'hFFFE;
        rom[70][10] = 16'h0011;
        rom[70][11] = 16'h0006;
        rom[70][12] = 16'h0024;
        rom[70][13] = 16'h0011;
        rom[70][14] = 16'h0011;
        rom[70][15] = 16'h0012;
        rom[70][16] = 16'hFFFC;
        rom[70][17] = 16'h0002;
        rom[70][18] = 16'h0016;
        rom[70][19] = 16'h0009;
        rom[70][20] = 16'h0029;
        rom[70][21] = 16'h000D;
        rom[70][22] = 16'hFFEC;
        rom[70][23] = 16'hFFDF;
        rom[70][24] = 16'hFFE1;
        rom[70][25] = 16'h0006;
        rom[70][26] = 16'h0003;
        rom[70][27] = 16'hFFEC;
        rom[70][28] = 16'hFFD1;
        rom[70][29] = 16'hFFE3;
        rom[70][30] = 16'h0029;
        rom[70][31] = 16'hFFD4;
        rom[70][32] = 16'h0006;
        rom[70][33] = 16'hFFF4;
        rom[70][34] = 16'h000C;
        rom[70][35] = 16'hFFD3;
        rom[70][36] = 16'h002E;
        rom[70][37] = 16'hFFEC;
        rom[70][38] = 16'h000F;
        rom[70][39] = 16'h002F;
        rom[70][40] = 16'hFFD7;
        rom[70][41] = 16'hFFF1;
        rom[70][42] = 16'hFFFB;
        rom[70][43] = 16'h0010;
        rom[70][44] = 16'h000D;
        rom[70][45] = 16'hFFCB;
        rom[70][46] = 16'h000E;
        rom[70][47] = 16'hFFDB;
        rom[70][48] = 16'h0004;
        rom[70][49] = 16'hFFE1;
        rom[70][50] = 16'h0015;
        rom[70][51] = 16'h0060;
        rom[70][52] = 16'h0006;
        rom[70][53] = 16'hFFFE;
        rom[70][54] = 16'hFFD6;
        rom[70][55] = 16'h000B;
        rom[70][56] = 16'hFFE8;
        rom[70][57] = 16'h002D;
        rom[70][58] = 16'hFFD0;
        rom[70][59] = 16'hFFF9;
        rom[70][60] = 16'h0030;
        rom[70][61] = 16'h0002;
        rom[70][62] = 16'hFFDC;
        rom[70][63] = 16'hFFD3;
        rom[70][64] = 16'hFFF1;
        rom[70][65] = 16'hFFFB;
        rom[70][66] = 16'h0003;
        rom[70][67] = 16'hFFFC;
        rom[70][68] = 16'h0017;
        rom[70][69] = 16'hFFDF;
        rom[70][70] = 16'hFFF4;
        rom[70][71] = 16'h0002;
        rom[70][72] = 16'hFFDF;
        rom[70][73] = 16'hFFE2;
        rom[70][74] = 16'hFFE8;
        rom[70][75] = 16'hFFE2;
        rom[70][76] = 16'h0008;
        rom[70][77] = 16'h000A;
        rom[70][78] = 16'h001F;
        rom[70][79] = 16'h0022;
        rom[70][80] = 16'hFFDA;
        rom[70][81] = 16'hFFE4;
        rom[70][82] = 16'hFFE5;
        rom[70][83] = 16'h000D;
        rom[70][84] = 16'h0029;
        rom[70][85] = 16'h0005;
        rom[70][86] = 16'hFFE5;
        rom[70][87] = 16'h000E;
        rom[70][88] = 16'h0010;
        rom[70][89] = 16'hFFE0;
        rom[70][90] = 16'hFFF4;
        rom[70][91] = 16'h0038;
        rom[70][92] = 16'hFFDE;
        rom[70][93] = 16'hFFBA;
        rom[70][94] = 16'h001F;
        rom[70][95] = 16'h001F;
        rom[70][96] = 16'h0003;
        rom[70][97] = 16'hFFA7;
        rom[70][98] = 16'hFFE5;
        rom[70][99] = 16'h001E;
        rom[70][100] = 16'hFFCE;
        rom[70][101] = 16'h0011;
        rom[70][102] = 16'hFFD0;
        rom[70][103] = 16'h0007;
        rom[70][104] = 16'h0028;
        rom[70][105] = 16'hFFC3;
        rom[70][106] = 16'hFFFE;
        rom[70][107] = 16'hFFFE;
        rom[70][108] = 16'hFFF1;
        rom[70][109] = 16'hFFF6;
        rom[70][110] = 16'hFFDB;
        rom[70][111] = 16'hFFE6;
        rom[70][112] = 16'h0023;
        rom[70][113] = 16'h002A;
        rom[70][114] = 16'hFFEC;
        rom[70][115] = 16'h0017;
        rom[70][116] = 16'h0002;
        rom[70][117] = 16'hFFDC;
        rom[70][118] = 16'h0005;
        rom[70][119] = 16'hFFC7;
        rom[70][120] = 16'h003C;
        rom[70][121] = 16'hFFD6;
        rom[70][122] = 16'hFFFC;
        rom[70][123] = 16'h0019;
        rom[70][124] = 16'hFFEA;
        rom[70][125] = 16'h001F;
        rom[70][126] = 16'hFFFE;
        rom[70][127] = 16'h0011;
        rom[71][0] = 16'hFFFE;
        rom[71][1] = 16'h0016;
        rom[71][2] = 16'hFFEC;
        rom[71][3] = 16'hFFF4;
        rom[71][4] = 16'hFFE1;
        rom[71][5] = 16'h0009;
        rom[71][6] = 16'h0001;
        rom[71][7] = 16'h0009;
        rom[71][8] = 16'h000C;
        rom[71][9] = 16'h001A;
        rom[71][10] = 16'hFFFA;
        rom[71][11] = 16'h001F;
        rom[71][12] = 16'hFFCD;
        rom[71][13] = 16'h000B;
        rom[71][14] = 16'h0008;
        rom[71][15] = 16'hFFE2;
        rom[71][16] = 16'hFFED;
        rom[71][17] = 16'hFFDF;
        rom[71][18] = 16'h0031;
        rom[71][19] = 16'hFFED;
        rom[71][20] = 16'h0012;
        rom[71][21] = 16'hFFEC;
        rom[71][22] = 16'h0038;
        rom[71][23] = 16'hFFAB;
        rom[71][24] = 16'hFFBE;
        rom[71][25] = 16'hFFFC;
        rom[71][26] = 16'h0001;
        rom[71][27] = 16'hFFD3;
        rom[71][28] = 16'h000A;
        rom[71][29] = 16'hFFE2;
        rom[71][30] = 16'hFFE9;
        rom[71][31] = 16'h000D;
        rom[71][32] = 16'h0027;
        rom[71][33] = 16'hFFDC;
        rom[71][34] = 16'hFFD7;
        rom[71][35] = 16'hFFF7;
        rom[71][36] = 16'h0005;
        rom[71][37] = 16'hFFC0;
        rom[71][38] = 16'h0005;
        rom[71][39] = 16'hFFDF;
        rom[71][40] = 16'hFFF6;
        rom[71][41] = 16'h0001;
        rom[71][42] = 16'h0026;
        rom[71][43] = 16'h000A;
        rom[71][44] = 16'hFFDA;
        rom[71][45] = 16'h0013;
        rom[71][46] = 16'hFFF1;
        rom[71][47] = 16'h0009;
        rom[71][48] = 16'hFFD8;
        rom[71][49] = 16'hFFF5;
        rom[71][50] = 16'hFFD9;
        rom[71][51] = 16'h001D;
        rom[71][52] = 16'h002E;
        rom[71][53] = 16'hFFF4;
        rom[71][54] = 16'h000D;
        rom[71][55] = 16'h0021;
        rom[71][56] = 16'hFFEA;
        rom[71][57] = 16'hFFEF;
        rom[71][58] = 16'h000A;
        rom[71][59] = 16'h0011;
        rom[71][60] = 16'hFFD7;
        rom[71][61] = 16'hFFC8;
        rom[71][62] = 16'hFFFA;
        rom[71][63] = 16'hFFE8;
        rom[71][64] = 16'hFFDF;
        rom[71][65] = 16'h0001;
        rom[71][66] = 16'h0019;
        rom[71][67] = 16'h0002;
        rom[71][68] = 16'hFFF3;
        rom[71][69] = 16'h0010;
        rom[71][70] = 16'hFFE4;
        rom[71][71] = 16'h0028;
        rom[71][72] = 16'hFFEA;
        rom[71][73] = 16'h000F;
        rom[71][74] = 16'h0021;
        rom[71][75] = 16'hFFBA;
        rom[71][76] = 16'hFFC4;
        rom[71][77] = 16'h001C;
        rom[71][78] = 16'h002B;
        rom[71][79] = 16'h000A;
        rom[71][80] = 16'h0033;
        rom[71][81] = 16'h0007;
        rom[71][82] = 16'hFFF6;
        rom[71][83] = 16'hFFF8;
        rom[71][84] = 16'h001A;
        rom[71][85] = 16'hFFFE;
        rom[71][86] = 16'h0022;
        rom[71][87] = 16'hFFFF;
        rom[71][88] = 16'hFFCD;
        rom[71][89] = 16'h0019;
        rom[71][90] = 16'hFFDC;
        rom[71][91] = 16'h0027;
        rom[71][92] = 16'hFFCE;
        rom[71][93] = 16'hFFF4;
        rom[71][94] = 16'hFFF7;
        rom[71][95] = 16'h003D;
        rom[71][96] = 16'h0026;
        rom[71][97] = 16'hFFFE;
        rom[71][98] = 16'hFFFE;
        rom[71][99] = 16'h0019;
        rom[71][100] = 16'h0027;
        rom[71][101] = 16'h001C;
        rom[71][102] = 16'hFFA8;
        rom[71][103] = 16'h0017;
        rom[71][104] = 16'h0014;
        rom[71][105] = 16'hFFB7;
        rom[71][106] = 16'hFFAF;
        rom[71][107] = 16'h0016;
        rom[71][108] = 16'hFFE0;
        rom[71][109] = 16'h000D;
        rom[71][110] = 16'hFFBD;
        rom[71][111] = 16'h001F;
        rom[71][112] = 16'h000C;
        rom[71][113] = 16'hFFFB;
        rom[71][114] = 16'hFFBD;
        rom[71][115] = 16'h0011;
        rom[71][116] = 16'hFFD7;
        rom[71][117] = 16'hFFD8;
        rom[71][118] = 16'hFFCD;
        rom[71][119] = 16'hFFD3;
        rom[71][120] = 16'hFFEF;
        rom[71][121] = 16'hFFD4;
        rom[71][122] = 16'h0017;
        rom[71][123] = 16'hFFBF;
        rom[71][124] = 16'h0007;
        rom[71][125] = 16'h0049;
        rom[71][126] = 16'hFFF4;
        rom[71][127] = 16'h0001;
        rom[72][0] = 16'hFFF9;
        rom[72][1] = 16'hFFD3;
        rom[72][2] = 16'h0023;
        rom[72][3] = 16'hFFFF;
        rom[72][4] = 16'h0010;
        rom[72][5] = 16'h0016;
        rom[72][6] = 16'hFFF4;
        rom[72][7] = 16'hFFB3;
        rom[72][8] = 16'h0009;
        rom[72][9] = 16'h0000;
        rom[72][10] = 16'h0006;
        rom[72][11] = 16'hFFDC;
        rom[72][12] = 16'hFFEE;
        rom[72][13] = 16'hFFC3;
        rom[72][14] = 16'hFFEF;
        rom[72][15] = 16'h0016;
        rom[72][16] = 16'h0007;
        rom[72][17] = 16'hFFB5;
        rom[72][18] = 16'hFF96;
        rom[72][19] = 16'hFFF2;
        rom[72][20] = 16'hFFE5;
        rom[72][21] = 16'hFFF7;
        rom[72][22] = 16'hFFE5;
        rom[72][23] = 16'hFFC7;
        rom[72][24] = 16'h000C;
        rom[72][25] = 16'h0007;
        rom[72][26] = 16'h0002;
        rom[72][27] = 16'h0007;
        rom[72][28] = 16'hFFE9;
        rom[72][29] = 16'h0017;
        rom[72][30] = 16'hFFD6;
        rom[72][31] = 16'h000A;
        rom[72][32] = 16'hFFD0;
        rom[72][33] = 16'hFFB8;
        rom[72][34] = 16'h000E;
        rom[72][35] = 16'hFFEA;
        rom[72][36] = 16'hFFD2;
        rom[72][37] = 16'hFFBC;
        rom[72][38] = 16'hFFB6;
        rom[72][39] = 16'h001E;
        rom[72][40] = 16'hFFF1;
        rom[72][41] = 16'h000A;
        rom[72][42] = 16'hFFF5;
        rom[72][43] = 16'hFFFC;
        rom[72][44] = 16'h0016;
        rom[72][45] = 16'h000B;
        rom[72][46] = 16'hFFCC;
        rom[72][47] = 16'h001F;
        rom[72][48] = 16'hFFDC;
        rom[72][49] = 16'hFFF6;
        rom[72][50] = 16'h0047;
        rom[72][51] = 16'hFFEB;
        rom[72][52] = 16'h0011;
        rom[72][53] = 16'h0000;
        rom[72][54] = 16'h0007;
        rom[72][55] = 16'h002C;
        rom[72][56] = 16'h000D;
        rom[72][57] = 16'h0022;
        rom[72][58] = 16'h0001;
        rom[72][59] = 16'hFFC9;
        rom[72][60] = 16'hFFEF;
        rom[72][61] = 16'h0011;
        rom[72][62] = 16'h0007;
        rom[72][63] = 16'hFFEA;
        rom[72][64] = 16'h0002;
        rom[72][65] = 16'hFFCD;
        rom[72][66] = 16'h003A;
        rom[72][67] = 16'h0017;
        rom[72][68] = 16'hFFFD;
        rom[72][69] = 16'h0002;
        rom[72][70] = 16'hFFEA;
        rom[72][71] = 16'hFFFE;
        rom[72][72] = 16'hFFE1;
        rom[72][73] = 16'h0009;
        rom[72][74] = 16'hFFDF;
        rom[72][75] = 16'hFFBC;
        rom[72][76] = 16'hFFCE;
        rom[72][77] = 16'hFFED;
        rom[72][78] = 16'h000D;
        rom[72][79] = 16'h0008;
        rom[72][80] = 16'hFFE7;
        rom[72][81] = 16'hFFF8;
        rom[72][82] = 16'hFFEF;
        rom[72][83] = 16'h0026;
        rom[72][84] = 16'hFFC8;
        rom[72][85] = 16'hFFF3;
        rom[72][86] = 16'h0006;
        rom[72][87] = 16'h0007;
        rom[72][88] = 16'hFFE5;
        rom[72][89] = 16'h0011;
        rom[72][90] = 16'hFFD1;
        rom[72][91] = 16'hFFEF;
        rom[72][92] = 16'hFFDF;
        rom[72][93] = 16'h000E;
        rom[72][94] = 16'hFFBC;
        rom[72][95] = 16'hFFF7;
        rom[72][96] = 16'hFFF4;
        rom[72][97] = 16'hFFF4;
        rom[72][98] = 16'h0002;
        rom[72][99] = 16'hFFD7;
        rom[72][100] = 16'hFFF0;
        rom[72][101] = 16'hFFF8;
        rom[72][102] = 16'hFFEA;
        rom[72][103] = 16'h0024;
        rom[72][104] = 16'hFFEB;
        rom[72][105] = 16'h001B;
        rom[72][106] = 16'hFFE5;
        rom[72][107] = 16'h0002;
        rom[72][108] = 16'hFFEA;
        rom[72][109] = 16'hFFEC;
        rom[72][110] = 16'hFFE8;
        rom[72][111] = 16'h0011;
        rom[72][112] = 16'hFFD9;
        rom[72][113] = 16'h0004;
        rom[72][114] = 16'hFFF1;
        rom[72][115] = 16'hFFF8;
        rom[72][116] = 16'hFFC7;
        rom[72][117] = 16'hFFE5;
        rom[72][118] = 16'hFFD9;
        rom[72][119] = 16'hFFFF;
        rom[72][120] = 16'hFFF0;
        rom[72][121] = 16'h000A;
        rom[72][122] = 16'hFFEE;
        rom[72][123] = 16'hFFDC;
        rom[72][124] = 16'hFFF5;
        rom[72][125] = 16'h0006;
        rom[72][126] = 16'h001A;
        rom[72][127] = 16'hFFFE;
        rom[73][0] = 16'hFFFC;
        rom[73][1] = 16'hFFF4;
        rom[73][2] = 16'h0004;
        rom[73][3] = 16'h0014;
        rom[73][4] = 16'hFFFE;
        rom[73][5] = 16'hFFC2;
        rom[73][6] = 16'h0014;
        rom[73][7] = 16'h0009;
        rom[73][8] = 16'hFFF2;
        rom[73][9] = 16'h0037;
        rom[73][10] = 16'h0025;
        rom[73][11] = 16'hFFC8;
        rom[73][12] = 16'hFFF6;
        rom[73][13] = 16'h000A;
        rom[73][14] = 16'hFFEF;
        rom[73][15] = 16'hFFD9;
        rom[73][16] = 16'h0033;
        rom[73][17] = 16'h0002;
        rom[73][18] = 16'h0022;
        rom[73][19] = 16'hFFFF;
        rom[73][20] = 16'hFFFD;
        rom[73][21] = 16'hFFEB;
        rom[73][22] = 16'hFFEA;
        rom[73][23] = 16'h0011;
        rom[73][24] = 16'hFFEA;
        rom[73][25] = 16'h000A;
        rom[73][26] = 16'hFFC8;
        rom[73][27] = 16'h0007;
        rom[73][28] = 16'hFFED;
        rom[73][29] = 16'h000A;
        rom[73][30] = 16'h002B;
        rom[73][31] = 16'h000C;
        rom[73][32] = 16'h0022;
        rom[73][33] = 16'hFFB5;
        rom[73][34] = 16'h0017;
        rom[73][35] = 16'hFFFB;
        rom[73][36] = 16'h002C;
        rom[73][37] = 16'hFFB1;
        rom[73][38] = 16'hFFD7;
        rom[73][39] = 16'h0016;
        rom[73][40] = 16'h0037;
        rom[73][41] = 16'hFFE8;
        rom[73][42] = 16'h0011;
        rom[73][43] = 16'hFFEB;
        rom[73][44] = 16'h0037;
        rom[73][45] = 16'h0017;
        rom[73][46] = 16'h0006;
        rom[73][47] = 16'hFFEF;
        rom[73][48] = 16'hFFF2;
        rom[73][49] = 16'h0014;
        rom[73][50] = 16'h0007;
        rom[73][51] = 16'h001B;
        rom[73][52] = 16'hFFE2;
        rom[73][53] = 16'h000C;
        rom[73][54] = 16'hFFEF;
        rom[73][55] = 16'h0001;
        rom[73][56] = 16'hFFE6;
        rom[73][57] = 16'hFFF4;
        rom[73][58] = 16'hFFB7;
        rom[73][59] = 16'h0012;
        rom[73][60] = 16'h0009;
        rom[73][61] = 16'h001A;
        rom[73][62] = 16'hFFFA;
        rom[73][63] = 16'h0006;
        rom[73][64] = 16'hFFFD;
        rom[73][65] = 16'h000F;
        rom[73][66] = 16'hFFC8;
        rom[73][67] = 16'hFFC1;
        rom[73][68] = 16'hFFDA;
        rom[73][69] = 16'hFFC4;
        rom[73][70] = 16'hFFF0;
        rom[73][71] = 16'hFFF0;
        rom[73][72] = 16'h0014;
        rom[73][73] = 16'hFFDE;
        rom[73][74] = 16'hFFDE;
        rom[73][75] = 16'hFFBB;
        rom[73][76] = 16'hFFEE;
        rom[73][77] = 16'h0010;
        rom[73][78] = 16'h0009;
        rom[73][79] = 16'hFFF4;
        rom[73][80] = 16'hFFE6;
        rom[73][81] = 16'hFFF0;
        rom[73][82] = 16'hFFCD;
        rom[73][83] = 16'h0015;
        rom[73][84] = 16'hFFE2;
        rom[73][85] = 16'h000D;
        rom[73][86] = 16'hFFEF;
        rom[73][87] = 16'hFFF6;
        rom[73][88] = 16'h001F;
        rom[73][89] = 16'hFFE1;
        rom[73][90] = 16'hFFF2;
        rom[73][91] = 16'h0024;
        rom[73][92] = 16'hFFE4;
        rom[73][93] = 16'hFFEF;
        rom[73][94] = 16'hFFF4;
        rom[73][95] = 16'hFFDB;
        rom[73][96] = 16'hFFED;
        rom[73][97] = 16'hFFE9;
        rom[73][98] = 16'h0014;
        rom[73][99] = 16'h0012;
        rom[73][100] = 16'hFFF4;
        rom[73][101] = 16'h000C;
        rom[73][102] = 16'h0024;
        rom[73][103] = 16'h0016;
        rom[73][104] = 16'h0001;
        rom[73][105] = 16'hFFEB;
        rom[73][106] = 16'hFFFF;
        rom[73][107] = 16'hFFD1;
        rom[73][108] = 16'hFFEB;
        rom[73][109] = 16'h0005;
        rom[73][110] = 16'hFFED;
        rom[73][111] = 16'hFFF2;
        rom[73][112] = 16'hFFD7;
        rom[73][113] = 16'hFFF5;
        rom[73][114] = 16'h0029;
        rom[73][115] = 16'h001B;
        rom[73][116] = 16'hFFB7;
        rom[73][117] = 16'hFFF3;
        rom[73][118] = 16'hFFB3;
        rom[73][119] = 16'hFFC7;
        rom[73][120] = 16'hFFFE;
        rom[73][121] = 16'hFFEC;
        rom[73][122] = 16'hFFFA;
        rom[73][123] = 16'hFFEF;
        rom[73][124] = 16'hFFE8;
        rom[73][125] = 16'hFFE2;
        rom[73][126] = 16'h0001;
        rom[73][127] = 16'h0032;
        rom[74][0] = 16'h0007;
        rom[74][1] = 16'hFFF2;
        rom[74][2] = 16'h002E;
        rom[74][3] = 16'hFFF9;
        rom[74][4] = 16'hFFFD;
        rom[74][5] = 16'h001D;
        rom[74][6] = 16'h0013;
        rom[74][7] = 16'hFFDA;
        rom[74][8] = 16'hFFF3;
        rom[74][9] = 16'h0027;
        rom[74][10] = 16'hFFC4;
        rom[74][11] = 16'hFFE0;
        rom[74][12] = 16'hFFD3;
        rom[74][13] = 16'h0002;
        rom[74][14] = 16'h0016;
        rom[74][15] = 16'h0024;
        rom[74][16] = 16'hFFF5;
        rom[74][17] = 16'hFFF2;
        rom[74][18] = 16'h0016;
        rom[74][19] = 16'h0026;
        rom[74][20] = 16'hFFC3;
        rom[74][21] = 16'h0016;
        rom[74][22] = 16'hFFFF;
        rom[74][23] = 16'hFFDE;
        rom[74][24] = 16'h000C;
        rom[74][25] = 16'h0016;
        rom[74][26] = 16'hFFFD;
        rom[74][27] = 16'hFFFE;
        rom[74][28] = 16'h0006;
        rom[74][29] = 16'h001A;
        rom[74][30] = 16'hFFF6;
        rom[74][31] = 16'hFFDE;
        rom[74][32] = 16'h0016;
        rom[74][33] = 16'hFFEC;
        rom[74][34] = 16'h0008;
        rom[74][35] = 16'hFFF5;
        rom[74][36] = 16'hFFD2;
        rom[74][37] = 16'h0027;
        rom[74][38] = 16'h0020;
        rom[74][39] = 16'h002B;
        rom[74][40] = 16'h000E;
        rom[74][41] = 16'hFFFA;
        rom[74][42] = 16'hFFDC;
        rom[74][43] = 16'hFFB8;
        rom[74][44] = 16'hFFF4;
        rom[74][45] = 16'h0016;
        rom[74][46] = 16'hFFEB;
        rom[74][47] = 16'h000A;
        rom[74][48] = 16'h0007;
        rom[74][49] = 16'hFFF5;
        rom[74][50] = 16'h002C;
        rom[74][51] = 16'hFFD7;
        rom[74][52] = 16'h0003;
        rom[74][53] = 16'h0033;
        rom[74][54] = 16'hFFD0;
        rom[74][55] = 16'h000C;
        rom[74][56] = 16'h0026;
        rom[74][57] = 16'hFFF4;
        rom[74][58] = 16'hFFD0;
        rom[74][59] = 16'hFFDC;
        rom[74][60] = 16'h0008;
        rom[74][61] = 16'hFFF3;
        rom[74][62] = 16'h0012;
        rom[74][63] = 16'hFFFA;
        rom[74][64] = 16'h0017;
        rom[74][65] = 16'hFFF6;
        rom[74][66] = 16'h0001;
        rom[74][67] = 16'h0007;
        rom[74][68] = 16'hFFDA;
        rom[74][69] = 16'h0011;
        rom[74][70] = 16'hFFF4;
        rom[74][71] = 16'h001B;
        rom[74][72] = 16'hFFDD;
        rom[74][73] = 16'h0010;
        rom[74][74] = 16'hFFF3;
        rom[74][75] = 16'h000B;
        rom[74][76] = 16'h0018;
        rom[74][77] = 16'hFFF9;
        rom[74][78] = 16'h0033;
        rom[74][79] = 16'hFFFB;
        rom[74][80] = 16'h0010;
        rom[74][81] = 16'hFFAD;
        rom[74][82] = 16'h000D;
        rom[74][83] = 16'hFFEF;
        rom[74][84] = 16'hFFEA;
        rom[74][85] = 16'h0017;
        rom[74][86] = 16'h0020;
        rom[74][87] = 16'hFFE6;
        rom[74][88] = 16'h0003;
        rom[74][89] = 16'h0008;
        rom[74][90] = 16'hFFF1;
        rom[74][91] = 16'h0002;
        rom[74][92] = 16'hFFF6;
        rom[74][93] = 16'hFFCC;
        rom[74][94] = 16'hFFD9;
        rom[74][95] = 16'hFFD6;
        rom[74][96] = 16'hFFC3;
        rom[74][97] = 16'hFFA9;
        rom[74][98] = 16'hFFDC;
        rom[74][99] = 16'h0069;
        rom[74][100] = 16'h0019;
        rom[74][101] = 16'h0018;
        rom[74][102] = 16'hFFEE;
        rom[74][103] = 16'hFFD8;
        rom[74][104] = 16'hFFEA;
        rom[74][105] = 16'h001E;
        rom[74][106] = 16'h001B;
        rom[74][107] = 16'hFFED;
        rom[74][108] = 16'hFFE5;
        rom[74][109] = 16'h0017;
        rom[74][110] = 16'h0000;
        rom[74][111] = 16'h0001;
        rom[74][112] = 16'h000E;
        rom[74][113] = 16'hFFF9;
        rom[74][114] = 16'hFFD7;
        rom[74][115] = 16'hFFD9;
        rom[74][116] = 16'hFFCF;
        rom[74][117] = 16'h0034;
        rom[74][118] = 16'h0025;
        rom[74][119] = 16'h0007;
        rom[74][120] = 16'h0010;
        rom[74][121] = 16'h000D;
        rom[74][122] = 16'h000A;
        rom[74][123] = 16'hFFDC;
        rom[74][124] = 16'hFFFF;
        rom[74][125] = 16'hFFF5;
        rom[74][126] = 16'h000F;
        rom[74][127] = 16'hFFF8;
        rom[75][0] = 16'hFFD4;
        rom[75][1] = 16'hFFCD;
        rom[75][2] = 16'hFFEB;
        rom[75][3] = 16'hFFC1;
        rom[75][4] = 16'h0014;
        rom[75][5] = 16'hFFF3;
        rom[75][6] = 16'hFFFB;
        rom[75][7] = 16'hFFF3;
        rom[75][8] = 16'hFFC9;
        rom[75][9] = 16'hFFDF;
        rom[75][10] = 16'hFFEF;
        rom[75][11] = 16'hFFFD;
        rom[75][12] = 16'hFFFA;
        rom[75][13] = 16'hFFF8;
        rom[75][14] = 16'h000C;
        rom[75][15] = 16'hFFE8;
        rom[75][16] = 16'hFFF4;
        rom[75][17] = 16'hFFDA;
        rom[75][18] = 16'h0035;
        rom[75][19] = 16'hFFAB;
        rom[75][20] = 16'h0032;
        rom[75][21] = 16'h000B;
        rom[75][22] = 16'hFFCD;
        rom[75][23] = 16'hFFD1;
        rom[75][24] = 16'hFFEB;
        rom[75][25] = 16'h0038;
        rom[75][26] = 16'hFFF9;
        rom[75][27] = 16'h0010;
        rom[75][28] = 16'hFFCC;
        rom[75][29] = 16'hFFCB;
        rom[75][30] = 16'h0046;
        rom[75][31] = 16'h001F;
        rom[75][32] = 16'hFFFF;
        rom[75][33] = 16'hFFF8;
        rom[75][34] = 16'hFFFD;
        rom[75][35] = 16'h0012;
        rom[75][36] = 16'hFFF4;
        rom[75][37] = 16'h000A;
        rom[75][38] = 16'hFFF6;
        rom[75][39] = 16'hFFF8;
        rom[75][40] = 16'hFFF4;
        rom[75][41] = 16'hFFDF;
        rom[75][42] = 16'hFFFA;
        rom[75][43] = 16'h0021;
        rom[75][44] = 16'h0029;
        rom[75][45] = 16'h0023;
        rom[75][46] = 16'hFFE6;
        rom[75][47] = 16'h000B;
        rom[75][48] = 16'h0007;
        rom[75][49] = 16'h0009;
        rom[75][50] = 16'hFFC4;
        rom[75][51] = 16'h0011;
        rom[75][52] = 16'hFFCD;
        rom[75][53] = 16'hFFD9;
        rom[75][54] = 16'h0004;
        rom[75][55] = 16'h0023;
        rom[75][56] = 16'h0026;
        rom[75][57] = 16'hFFF7;
        rom[75][58] = 16'h0028;
        rom[75][59] = 16'h0032;
        rom[75][60] = 16'h0033;
        rom[75][61] = 16'hFFFE;
        rom[75][62] = 16'hFFD8;
        rom[75][63] = 16'hFFEE;
        rom[75][64] = 16'hFFE1;
        rom[75][65] = 16'hFFE9;
        rom[75][66] = 16'h0002;
        rom[75][67] = 16'h000B;
        rom[75][68] = 16'hFFB5;
        rom[75][69] = 16'hFFFE;
        rom[75][70] = 16'hFFE1;
        rom[75][71] = 16'hFFD5;
        rom[75][72] = 16'h002B;
        rom[75][73] = 16'h0012;
        rom[75][74] = 16'hFFB5;
        rom[75][75] = 16'hFFFE;
        rom[75][76] = 16'hFFE2;
        rom[75][77] = 16'h0011;
        rom[75][78] = 16'hFFF4;
        rom[75][79] = 16'h001F;
        rom[75][80] = 16'hFFC0;
        rom[75][81] = 16'hFFF1;
        rom[75][82] = 16'h0002;
        rom[75][83] = 16'h0022;
        rom[75][84] = 16'h0000;
        rom[75][85] = 16'h000F;
        rom[75][86] = 16'hFFED;
        rom[75][87] = 16'hFFD3;
        rom[75][88] = 16'h004C;
        rom[75][89] = 16'hFFDE;
        rom[75][90] = 16'h0010;
        rom[75][91] = 16'hFFAF;
        rom[75][92] = 16'h001A;
        rom[75][93] = 16'hFFC8;
        rom[75][94] = 16'hFFF4;
        rom[75][95] = 16'hFFE3;
        rom[75][96] = 16'hFFC7;
        rom[75][97] = 16'hFFB3;
        rom[75][98] = 16'hFFF0;
        rom[75][99] = 16'h0002;
        rom[75][100] = 16'hFFF0;
        rom[75][101] = 16'hFFDC;
        rom[75][102] = 16'hFFF6;
        rom[75][103] = 16'hFFE1;
        rom[75][104] = 16'hFFE9;
        rom[75][105] = 16'hFF99;
        rom[75][106] = 16'hFFD3;
        rom[75][107] = 16'h0005;
        rom[75][108] = 16'hFFFD;
        rom[75][109] = 16'h0021;
        rom[75][110] = 16'hFFE5;
        rom[75][111] = 16'hFFE7;
        rom[75][112] = 16'h000C;
        rom[75][113] = 16'h0001;
        rom[75][114] = 16'h0012;
        rom[75][115] = 16'h0015;
        rom[75][116] = 16'hFFE8;
        rom[75][117] = 16'hFFFA;
        rom[75][118] = 16'hFFFC;
        rom[75][119] = 16'hFFEE;
        rom[75][120] = 16'h003D;
        rom[75][121] = 16'hFFB5;
        rom[75][122] = 16'h0009;
        rom[75][123] = 16'h0011;
        rom[75][124] = 16'hFFE3;
        rom[75][125] = 16'hFFF9;
        rom[75][126] = 16'hFFE8;
        rom[75][127] = 16'h001C;
        rom[76][0] = 16'hFFDC;
        rom[76][1] = 16'h0005;
        rom[76][2] = 16'h0004;
        rom[76][3] = 16'h0009;
        rom[76][4] = 16'hFFE5;
        rom[76][5] = 16'hFFFD;
        rom[76][6] = 16'hFFCD;
        rom[76][7] = 16'hFFF2;
        rom[76][8] = 16'h0001;
        rom[76][9] = 16'h0012;
        rom[76][10] = 16'h0016;
        rom[76][11] = 16'hFFB4;
        rom[76][12] = 16'h000C;
        rom[76][13] = 16'hFFFC;
        rom[76][14] = 16'hFFD5;
        rom[76][15] = 16'h0007;
        rom[76][16] = 16'hFFBE;
        rom[76][17] = 16'h000D;
        rom[76][18] = 16'h0007;
        rom[76][19] = 16'h0002;
        rom[76][20] = 16'h0012;
        rom[76][21] = 16'hFFF6;
        rom[76][22] = 16'h0033;
        rom[76][23] = 16'hFFF9;
        rom[76][24] = 16'hFFDD;
        rom[76][25] = 16'h0000;
        rom[76][26] = 16'h0006;
        rom[76][27] = 16'hFFF1;
        rom[76][28] = 16'hFFF4;
        rom[76][29] = 16'h0015;
        rom[76][30] = 16'hFFD5;
        rom[76][31] = 16'hFFCA;
        rom[76][32] = 16'h002B;
        rom[76][33] = 16'hFFF7;
        rom[76][34] = 16'hFFE3;
        rom[76][35] = 16'h0025;
        rom[76][36] = 16'hFFDD;
        rom[76][37] = 16'hFFDD;
        rom[76][38] = 16'h0016;
        rom[76][39] = 16'hFFFE;
        rom[76][40] = 16'h001B;
        rom[76][41] = 16'h0033;
        rom[76][42] = 16'h001B;
        rom[76][43] = 16'h000E;
        rom[76][44] = 16'h0002;
        rom[76][45] = 16'h000F;
        rom[76][46] = 16'hFFFA;
        rom[76][47] = 16'h0038;
        rom[76][48] = 16'hFFE0;
        rom[76][49] = 16'hFFE8;
        rom[76][50] = 16'h0014;
        rom[76][51] = 16'hFFE4;
        rom[76][52] = 16'hFFD2;
        rom[76][53] = 16'hFFE6;
        rom[76][54] = 16'h002A;
        rom[76][55] = 16'h0024;
        rom[76][56] = 16'hFFC9;
        rom[76][57] = 16'hFFEA;
        rom[76][58] = 16'h000B;
        rom[76][59] = 16'hFFE1;
        rom[76][60] = 16'hFFB9;
        rom[76][61] = 16'hFFFE;
        rom[76][62] = 16'h0008;
        rom[76][63] = 16'hFFF8;
        rom[76][64] = 16'h0024;
        rom[76][65] = 16'hFFE0;
        rom[76][66] = 16'h0004;
        rom[76][67] = 16'h0010;
        rom[76][68] = 16'hFFD2;
        rom[76][69] = 16'hFFF9;
        rom[76][70] = 16'hFFEF;
        rom[76][71] = 16'h002B;
        rom[76][72] = 16'hFFB0;
        rom[76][73] = 16'h0019;
        rom[76][74] = 16'hFFDC;
        rom[76][75] = 16'h0014;
        rom[76][76] = 16'hFFEF;
        rom[76][77] = 16'hFFD9;
        rom[76][78] = 16'h001F;
        rom[76][79] = 16'h0002;
        rom[76][80] = 16'h002C;
        rom[76][81] = 16'hFFE1;
        rom[76][82] = 16'hFFF9;
        rom[76][83] = 16'h0026;
        rom[76][84] = 16'h000A;
        rom[76][85] = 16'hFFEB;
        rom[76][86] = 16'hFFF2;
        rom[76][87] = 16'hFFEF;
        rom[76][88] = 16'h0029;
        rom[76][89] = 16'h0014;
        rom[76][90] = 16'hFFFC;
        rom[76][91] = 16'hFFBC;
        rom[76][92] = 16'hFFF2;
        rom[76][93] = 16'h0026;
        rom[76][94] = 16'hFFDF;
        rom[76][95] = 16'hFFF4;
        rom[76][96] = 16'h004E;
        rom[76][97] = 16'hFFEA;
        rom[76][98] = 16'hFFCD;
        rom[76][99] = 16'hFFEF;
        rom[76][100] = 16'h000C;
        rom[76][101] = 16'h0004;
        rom[76][102] = 16'hFFF0;
        rom[76][103] = 16'hFFF0;
        rom[76][104] = 16'hFFE5;
        rom[76][105] = 16'hFFF4;
        rom[76][106] = 16'hFFEC;
        rom[76][107] = 16'hFFE3;
        rom[76][108] = 16'hFFD6;
        rom[76][109] = 16'h0014;
        rom[76][110] = 16'hFFE2;
        rom[76][111] = 16'hFFDD;
        rom[76][112] = 16'hFFEF;
        rom[76][113] = 16'h001B;
        rom[76][114] = 16'hFFED;
        rom[76][115] = 16'hFFF4;
        rom[76][116] = 16'h0008;
        rom[76][117] = 16'h0002;
        rom[76][118] = 16'h0032;
        rom[76][119] = 16'h0025;
        rom[76][120] = 16'hFFC7;
        rom[76][121] = 16'hFFD7;
        rom[76][122] = 16'hFFDB;
        rom[76][123] = 16'hFFD7;
        rom[76][124] = 16'hFFD5;
        rom[76][125] = 16'h0004;
        rom[76][126] = 16'h0020;
        rom[76][127] = 16'h000D;
        rom[77][0] = 16'hFFEE;
        rom[77][1] = 16'h0013;
        rom[77][2] = 16'h0003;
        rom[77][3] = 16'hFFF2;
        rom[77][4] = 16'hFFE9;
        rom[77][5] = 16'hFFE7;
        rom[77][6] = 16'h0004;
        rom[77][7] = 16'hFFE8;
        rom[77][8] = 16'h000D;
        rom[77][9] = 16'hFFC5;
        rom[77][10] = 16'h0016;
        rom[77][11] = 16'hFFF6;
        rom[77][12] = 16'hFFF3;
        rom[77][13] = 16'hFFD1;
        rom[77][14] = 16'h0017;
        rom[77][15] = 16'hFFED;
        rom[77][16] = 16'h0024;
        rom[77][17] = 16'hFFE5;
        rom[77][18] = 16'hFFF1;
        rom[77][19] = 16'h000C;
        rom[77][20] = 16'h002C;
        rom[77][21] = 16'h0003;
        rom[77][22] = 16'hFFDA;
        rom[77][23] = 16'hFFE7;
        rom[77][24] = 16'hFFFE;
        rom[77][25] = 16'h002A;
        rom[77][26] = 16'h0036;
        rom[77][27] = 16'h000F;
        rom[77][28] = 16'h0004;
        rom[77][29] = 16'h0002;
        rom[77][30] = 16'hFFFA;
        rom[77][31] = 16'h0013;
        rom[77][32] = 16'h0008;
        rom[77][33] = 16'hFFE8;
        rom[77][34] = 16'h0015;
        rom[77][35] = 16'hFFED;
        rom[77][36] = 16'h0014;
        rom[77][37] = 16'h003D;
        rom[77][38] = 16'hFFCC;
        rom[77][39] = 16'h0011;
        rom[77][40] = 16'h0002;
        rom[77][41] = 16'hFFEF;
        rom[77][42] = 16'h0007;
        rom[77][43] = 16'h0007;
        rom[77][44] = 16'h000E;
        rom[77][45] = 16'hFFE0;
        rom[77][46] = 16'hFFEB;
        rom[77][47] = 16'h0035;
        rom[77][48] = 16'hFFD0;
        rom[77][49] = 16'hFFCE;
        rom[77][50] = 16'hFFFE;
        rom[77][51] = 16'hFFF9;
        rom[77][52] = 16'h0010;
        rom[77][53] = 16'hFFFC;
        rom[77][54] = 16'hFFD2;
        rom[77][55] = 16'hFFF9;
        rom[77][56] = 16'hFFEC;
        rom[77][57] = 16'hFFEC;
        rom[77][58] = 16'hFFC8;
        rom[77][59] = 16'hFFFD;
        rom[77][60] = 16'hFFE6;
        rom[77][61] = 16'hFFEF;
        rom[77][62] = 16'h0026;
        rom[77][63] = 16'hFFD6;
        rom[77][64] = 16'hFFC8;
        rom[77][65] = 16'hFFF4;
        rom[77][66] = 16'hFFDB;
        rom[77][67] = 16'hFFE7;
        rom[77][68] = 16'hFFFB;
        rom[77][69] = 16'hFFFC;
        rom[77][70] = 16'hFFAB;
        rom[77][71] = 16'h000F;
        rom[77][72] = 16'h0001;
        rom[77][73] = 16'hFFCE;
        rom[77][74] = 16'h0005;
        rom[77][75] = 16'hFFF7;
        rom[77][76] = 16'hFFEC;
        rom[77][77] = 16'hFFE0;
        rom[77][78] = 16'h0021;
        rom[77][79] = 16'hFFDD;
        rom[77][80] = 16'h0024;
        rom[77][81] = 16'hFFCD;
        rom[77][82] = 16'h0019;
        rom[77][83] = 16'hFFF2;
        rom[77][84] = 16'hFFC7;
        rom[77][85] = 16'h0008;
        rom[77][86] = 16'h0006;
        rom[77][87] = 16'hFFF1;
        rom[77][88] = 16'h0012;
        rom[77][89] = 16'hFFE4;
        rom[77][90] = 16'h0009;
        rom[77][91] = 16'hFFFE;
        rom[77][92] = 16'h000E;
        rom[77][93] = 16'hFFF5;
        rom[77][94] = 16'h000B;
        rom[77][95] = 16'hFFFE;
        rom[77][96] = 16'h0006;
        rom[77][97] = 16'h0006;
        rom[77][98] = 16'h0029;
        rom[77][99] = 16'hFFDB;
        rom[77][100] = 16'h0019;
        rom[77][101] = 16'h0015;
        rom[77][102] = 16'hFFF4;
        rom[77][103] = 16'hFFD4;
        rom[77][104] = 16'hFFE0;
        rom[77][105] = 16'hFFE6;
        rom[77][106] = 16'hFFF3;
        rom[77][107] = 16'hFFEB;
        rom[77][108] = 16'h0004;
        rom[77][109] = 16'hFFEA;
        rom[77][110] = 16'hFFD9;
        rom[77][111] = 16'h0024;
        rom[77][112] = 16'h002B;
        rom[77][113] = 16'hFFD6;
        rom[77][114] = 16'h0005;
        rom[77][115] = 16'h0015;
        rom[77][116] = 16'hFFD6;
        rom[77][117] = 16'h0032;
        rom[77][118] = 16'hFFFA;
        rom[77][119] = 16'hFFF0;
        rom[77][120] = 16'hFFD4;
        rom[77][121] = 16'h000E;
        rom[77][122] = 16'hFFE3;
        rom[77][123] = 16'hFFFE;
        rom[77][124] = 16'hFFE3;
        rom[77][125] = 16'hFFCB;
        rom[77][126] = 16'h0011;
        rom[77][127] = 16'h0000;
        rom[78][0] = 16'hFFFC;
        rom[78][1] = 16'h0009;
        rom[78][2] = 16'hFFF0;
        rom[78][3] = 16'hFFF5;
        rom[78][4] = 16'h0003;
        rom[78][5] = 16'h0016;
        rom[78][6] = 16'hFFDE;
        rom[78][7] = 16'hFFDB;
        rom[78][8] = 16'hFFF8;
        rom[78][9] = 16'h0015;
        rom[78][10] = 16'hFFFD;
        rom[78][11] = 16'h000C;
        rom[78][12] = 16'hFFC5;
        rom[78][13] = 16'h0002;
        rom[78][14] = 16'h0016;
        rom[78][15] = 16'hFFCE;
        rom[78][16] = 16'hFFEA;
        rom[78][17] = 16'hFFFE;
        rom[78][18] = 16'hFFFB;
        rom[78][19] = 16'hFFFB;
        rom[78][20] = 16'hFFF9;
        rom[78][21] = 16'hFFEE;
        rom[78][22] = 16'hFFCD;
        rom[78][23] = 16'h0002;
        rom[78][24] = 16'h000C;
        rom[78][25] = 16'hFFFA;
        rom[78][26] = 16'h001D;
        rom[78][27] = 16'hFFB9;
        rom[78][28] = 16'h0037;
        rom[78][29] = 16'h0018;
        rom[78][30] = 16'hFFDC;
        rom[78][31] = 16'hFFD2;
        rom[78][32] = 16'h0015;
        rom[78][33] = 16'hFFF4;
        rom[78][34] = 16'hFFE2;
        rom[78][35] = 16'hFFD1;
        rom[78][36] = 16'hFFD6;
        rom[78][37] = 16'h0010;
        rom[78][38] = 16'hFFCE;
        rom[78][39] = 16'h0000;
        rom[78][40] = 16'h0016;
        rom[78][41] = 16'hFFE7;
        rom[78][42] = 16'h0013;
        rom[78][43] = 16'h0007;
        rom[78][44] = 16'h0002;
        rom[78][45] = 16'hFFFD;
        rom[78][46] = 16'hFFE9;
        rom[78][47] = 16'hFFEB;
        rom[78][48] = 16'hFFC8;
        rom[78][49] = 16'hFFFA;
        rom[78][50] = 16'hFFD2;
        rom[78][51] = 16'hFFF5;
        rom[78][52] = 16'h0001;
        rom[78][53] = 16'h000D;
        rom[78][54] = 16'hFFF9;
        rom[78][55] = 16'hFFD9;
        rom[78][56] = 16'hFFF4;
        rom[78][57] = 16'hFFE1;
        rom[78][58] = 16'hFFED;
        rom[78][59] = 16'h0002;
        rom[78][60] = 16'h0007;
        rom[78][61] = 16'hFFDC;
        rom[78][62] = 16'hFFF0;
        rom[78][63] = 16'hFFE0;
        rom[78][64] = 16'h0022;
        rom[78][65] = 16'hFFF9;
        rom[78][66] = 16'h0016;
        rom[78][67] = 16'h0010;
        rom[78][68] = 16'h0024;
        rom[78][69] = 16'h0012;
        rom[78][70] = 16'hFFDC;
        rom[78][71] = 16'hFFD7;
        rom[78][72] = 16'hFFE1;
        rom[78][73] = 16'hFFFF;
        rom[78][74] = 16'hFFFF;
        rom[78][75] = 16'h0012;
        rom[78][76] = 16'hFFFA;
        rom[78][77] = 16'h0014;
        rom[78][78] = 16'h0041;
        rom[78][79] = 16'h0003;
        rom[78][80] = 16'hFFEF;
        rom[78][81] = 16'h0001;
        rom[78][82] = 16'h0015;
        rom[78][83] = 16'h0006;
        rom[78][84] = 16'hFFE9;
        rom[78][85] = 16'hFFDA;
        rom[78][86] = 16'h0013;
        rom[78][87] = 16'hFFEB;
        rom[78][88] = 16'h0003;
        rom[78][89] = 16'hFFD2;
        rom[78][90] = 16'hFFFE;
        rom[78][91] = 16'hFFE5;
        rom[78][92] = 16'h0025;
        rom[78][93] = 16'hFFD0;
        rom[78][94] = 16'h0011;
        rom[78][95] = 16'hFFFF;
        rom[78][96] = 16'h0002;
        rom[78][97] = 16'hFFE5;
        rom[78][98] = 16'hFFB5;
        rom[78][99] = 16'hFFC9;
        rom[78][100] = 16'h000C;
        rom[78][101] = 16'hFFFB;
        rom[78][102] = 16'hFFD7;
        rom[78][103] = 16'h0010;
        rom[78][104] = 16'hFFEA;
        rom[78][105] = 16'hFFF5;
        rom[78][106] = 16'h0024;
        rom[78][107] = 16'hFFC7;
        rom[78][108] = 16'hFFC8;
        rom[78][109] = 16'hFFF9;
        rom[78][110] = 16'h0002;
        rom[78][111] = 16'hFFE9;
        rom[78][112] = 16'hFFE5;
        rom[78][113] = 16'hFFF5;
        rom[78][114] = 16'hFFF5;
        rom[78][115] = 16'hFFC9;
        rom[78][116] = 16'h000D;
        rom[78][117] = 16'h0020;
        rom[78][118] = 16'h0004;
        rom[78][119] = 16'hFFDC;
        rom[78][120] = 16'hFFEE;
        rom[78][121] = 16'hFFF5;
        rom[78][122] = 16'h000E;
        rom[78][123] = 16'hFFF9;
        rom[78][124] = 16'hFFDE;
        rom[78][125] = 16'hFFD5;
        rom[78][126] = 16'hFFE0;
        rom[78][127] = 16'hFFC1;
        rom[79][0] = 16'hFFC6;
        rom[79][1] = 16'hFFCE;
        rom[79][2] = 16'hFFF7;
        rom[79][3] = 16'hFFDA;
        rom[79][4] = 16'hFFF9;
        rom[79][5] = 16'h0015;
        rom[79][6] = 16'h000F;
        rom[79][7] = 16'h000B;
        rom[79][8] = 16'hFFE5;
        rom[79][9] = 16'h002A;
        rom[79][10] = 16'hFFDC;
        rom[79][11] = 16'hFFFD;
        rom[79][12] = 16'hFFFF;
        rom[79][13] = 16'h0016;
        rom[79][14] = 16'h0011;
        rom[79][15] = 16'hFFDC;
        rom[79][16] = 16'h001D;
        rom[79][17] = 16'hFFF6;
        rom[79][18] = 16'hFFE8;
        rom[79][19] = 16'hFFD7;
        rom[79][20] = 16'hFFF9;
        rom[79][21] = 16'hFFED;
        rom[79][22] = 16'hFFF4;
        rom[79][23] = 16'h0002;
        rom[79][24] = 16'h000F;
        rom[79][25] = 16'h0016;
        rom[79][26] = 16'hFFCA;
        rom[79][27] = 16'h001F;
        rom[79][28] = 16'h0033;
        rom[79][29] = 16'h0005;
        rom[79][30] = 16'h0002;
        rom[79][31] = 16'h0007;
        rom[79][32] = 16'h0003;
        rom[79][33] = 16'hFFF5;
        rom[79][34] = 16'h0007;
        rom[79][35] = 16'h0038;
        rom[79][36] = 16'h0002;
        rom[79][37] = 16'hFFD8;
        rom[79][38] = 16'h0048;
        rom[79][39] = 16'hFFFF;
        rom[79][40] = 16'h0017;
        rom[79][41] = 16'hFFEC;
        rom[79][42] = 16'hFFF4;
        rom[79][43] = 16'hFFEE;
        rom[79][44] = 16'h000C;
        rom[79][45] = 16'h0014;
        rom[79][46] = 16'h0007;
        rom[79][47] = 16'h0001;
        rom[79][48] = 16'h0041;
        rom[79][49] = 16'h0001;
        rom[79][50] = 16'h003D;
        rom[79][51] = 16'hFFEB;
        rom[79][52] = 16'h0002;
        rom[79][53] = 16'h000E;
        rom[79][54] = 16'h0014;
        rom[79][55] = 16'h0014;
        rom[79][56] = 16'hFFBB;
        rom[79][57] = 16'h000C;
        rom[79][58] = 16'h000A;
        rom[79][59] = 16'hFFE5;
        rom[79][60] = 16'hFFE0;
        rom[79][61] = 16'hFFF9;
        rom[79][62] = 16'h0008;
        rom[79][63] = 16'h0004;
        rom[79][64] = 16'hFFE5;
        rom[79][65] = 16'h0002;
        rom[79][66] = 16'hFFCD;
        rom[79][67] = 16'hFFCD;
        rom[79][68] = 16'hFFF3;
        rom[79][69] = 16'hFFAF;
        rom[79][70] = 16'h0006;
        rom[79][71] = 16'h0002;
        rom[79][72] = 16'hFFBF;
        rom[79][73] = 16'hFFEC;
        rom[79][74] = 16'h0000;
        rom[79][75] = 16'h000C;
        rom[79][76] = 16'hFFE0;
        rom[79][77] = 16'hFFFA;
        rom[79][78] = 16'hFFCA;
        rom[79][79] = 16'hFFF4;
        rom[79][80] = 16'hFFE3;
        rom[79][81] = 16'hFFEF;
        rom[79][82] = 16'hFFE3;
        rom[79][83] = 16'h0010;
        rom[79][84] = 16'hFFD0;
        rom[79][85] = 16'h0042;
        rom[79][86] = 16'h0013;
        rom[79][87] = 16'h0016;
        rom[79][88] = 16'hFFF4;
        rom[79][89] = 16'h0016;
        rom[79][90] = 16'hFFEE;
        rom[79][91] = 16'hFFF6;
        rom[79][92] = 16'h001B;
        rom[79][93] = 16'h000F;
        rom[79][94] = 16'hFFF5;
        rom[79][95] = 16'h001C;
        rom[79][96] = 16'hFFFC;
        rom[79][97] = 16'h0002;
        rom[79][98] = 16'hFFDB;
        rom[79][99] = 16'hFFB6;
        rom[79][100] = 16'h000C;
        rom[79][101] = 16'h000C;
        rom[79][102] = 16'h0025;
        rom[79][103] = 16'hFFEE;
        rom[79][104] = 16'hFFEA;
        rom[79][105] = 16'h0002;
        rom[79][106] = 16'h0011;
        rom[79][107] = 16'hFFE1;
        rom[79][108] = 16'h001A;
        rom[79][109] = 16'h0019;
        rom[79][110] = 16'h0009;
        rom[79][111] = 16'hFFCF;
        rom[79][112] = 16'h0027;
        rom[79][113] = 16'h0020;
        rom[79][114] = 16'h002E;
        rom[79][115] = 16'hFFFB;
        rom[79][116] = 16'h0017;
        rom[79][117] = 16'h000F;
        rom[79][118] = 16'h001C;
        rom[79][119] = 16'h001D;
        rom[79][120] = 16'h0014;
        rom[79][121] = 16'h0027;
        rom[79][122] = 16'hFFF9;
        rom[79][123] = 16'h003C;
        rom[79][124] = 16'h0003;
        rom[79][125] = 16'hFFF4;
        rom[79][126] = 16'h000B;
        rom[79][127] = 16'hFFD9;
        rom[80][0] = 16'hFFEC;
        rom[80][1] = 16'hFFCF;
        rom[80][2] = 16'hFFFB;
        rom[80][3] = 16'hFFFE;
        rom[80][4] = 16'h0006;
        rom[80][5] = 16'hFFFB;
        rom[80][6] = 16'h0016;
        rom[80][7] = 16'hFFB6;
        rom[80][8] = 16'hFFDC;
        rom[80][9] = 16'hFFE1;
        rom[80][10] = 16'h001E;
        rom[80][11] = 16'h0008;
        rom[80][12] = 16'h0027;
        rom[80][13] = 16'hFFBE;
        rom[80][14] = 16'hFFE1;
        rom[80][15] = 16'h0014;
        rom[80][16] = 16'h0029;
        rom[80][17] = 16'hFFCD;
        rom[80][18] = 16'hFFEA;
        rom[80][19] = 16'hFFF1;
        rom[80][20] = 16'hFFFB;
        rom[80][21] = 16'h0000;
        rom[80][22] = 16'hFFEB;
        rom[80][23] = 16'hFFEE;
        rom[80][24] = 16'h0005;
        rom[80][25] = 16'hFFEA;
        rom[80][26] = 16'hFFE8;
        rom[80][27] = 16'h0010;
        rom[80][28] = 16'hFFEF;
        rom[80][29] = 16'hFFA1;
        rom[80][30] = 16'h0012;
        rom[80][31] = 16'hFFE0;
        rom[80][32] = 16'hFFDC;
        rom[80][33] = 16'hFFDE;
        rom[80][34] = 16'hFFFC;
        rom[80][35] = 16'hFFEF;
        rom[80][36] = 16'hFFF7;
        rom[80][37] = 16'hFFDF;
        rom[80][38] = 16'hFFF7;
        rom[80][39] = 16'h002E;
        rom[80][40] = 16'hFFDD;
        rom[80][41] = 16'h000D;
        rom[80][42] = 16'h0006;
        rom[80][43] = 16'h000B;
        rom[80][44] = 16'h000D;
        rom[80][45] = 16'h000D;
        rom[80][46] = 16'h0008;
        rom[80][47] = 16'hFFFC;
        rom[80][48] = 16'hFFF1;
        rom[80][49] = 16'hFFB8;
        rom[80][50] = 16'h001B;
        rom[80][51] = 16'h0029;
        rom[80][52] = 16'h0006;
        rom[80][53] = 16'h0011;
        rom[80][54] = 16'h0016;
        rom[80][55] = 16'hFFEF;
        rom[80][56] = 16'h0008;
        rom[80][57] = 16'h0027;
        rom[80][58] = 16'h001B;
        rom[80][59] = 16'hFFFF;
        rom[80][60] = 16'h0022;
        rom[80][61] = 16'hFFF3;
        rom[80][62] = 16'hFFF0;
        rom[80][63] = 16'hFFC8;
        rom[80][64] = 16'h005B;
        rom[80][65] = 16'h0002;
        rom[80][66] = 16'hFFFD;
        rom[80][67] = 16'hFFFD;
        rom[80][68] = 16'hFFEF;
        rom[80][69] = 16'hFFE1;
        rom[80][70] = 16'hFFF2;
        rom[80][71] = 16'hFFF4;
        rom[80][72] = 16'h0004;
        rom[80][73] = 16'hFFEC;
        rom[80][74] = 16'hFFE1;
        rom[80][75] = 16'hFFF7;
        rom[80][76] = 16'h0016;
        rom[80][77] = 16'h0014;
        rom[80][78] = 16'h0036;
        rom[80][79] = 16'h0021;
        rom[80][80] = 16'hFFFC;
        rom[80][81] = 16'h000A;
        rom[80][82] = 16'hFFBA;
        rom[80][83] = 16'h0005;
        rom[80][84] = 16'h0028;
        rom[80][85] = 16'h000C;
        rom[80][86] = 16'hFFC3;
        rom[80][87] = 16'h001D;
        rom[80][88] = 16'hFFFD;
        rom[80][89] = 16'h002C;
        rom[80][90] = 16'hFFBA;
        rom[80][91] = 16'h001E;
        rom[80][92] = 16'h0027;
        rom[80][93] = 16'hFFBF;
        rom[80][94] = 16'hFFF1;
        rom[80][95] = 16'hFFDF;
        rom[80][96] = 16'h000E;
        rom[80][97] = 16'hFFE8;
        rom[80][98] = 16'hFFEF;
        rom[80][99] = 16'h0005;
        rom[80][100] = 16'hFFC3;
        rom[80][101] = 16'hFFD0;
        rom[80][102] = 16'hFFA6;
        rom[80][103] = 16'hFFCF;
        rom[80][104] = 16'h002B;
        rom[80][105] = 16'h000C;
        rom[80][106] = 16'hFFF4;
        rom[80][107] = 16'h0009;
        rom[80][108] = 16'hFFE4;
        rom[80][109] = 16'hFFD1;
        rom[80][110] = 16'hFFEF;
        rom[80][111] = 16'hFFE3;
        rom[80][112] = 16'h0007;
        rom[80][113] = 16'h002D;
        rom[80][114] = 16'hFFD3;
        rom[80][115] = 16'h000D;
        rom[80][116] = 16'hFFFF;
        rom[80][117] = 16'hFFDD;
        rom[80][118] = 16'h0014;
        rom[80][119] = 16'h0016;
        rom[80][120] = 16'h0029;
        rom[80][121] = 16'h0013;
        rom[80][122] = 16'h002A;
        rom[80][123] = 16'h000E;
        rom[80][124] = 16'h0016;
        rom[80][125] = 16'h001C;
        rom[80][126] = 16'h001E;
        rom[80][127] = 16'h001D;
        rom[81][0] = 16'h0024;
        rom[81][1] = 16'hFFBF;
        rom[81][2] = 16'hFFC8;
        rom[81][3] = 16'hFFDF;
        rom[81][4] = 16'hFFEF;
        rom[81][5] = 16'hFFED;
        rom[81][6] = 16'h0011;
        rom[81][7] = 16'hFFE4;
        rom[81][8] = 16'hFFD2;
        rom[81][9] = 16'hFFDD;
        rom[81][10] = 16'hFFED;
        rom[81][11] = 16'h000D;
        rom[81][12] = 16'h0005;
        rom[81][13] = 16'hFFE1;
        rom[81][14] = 16'h0022;
        rom[81][15] = 16'hFFE6;
        rom[81][16] = 16'hFFED;
        rom[81][17] = 16'hFFFE;
        rom[81][18] = 16'hFFF3;
        rom[81][19] = 16'hFFD3;
        rom[81][20] = 16'hFFFA;
        rom[81][21] = 16'hFFDC;
        rom[81][22] = 16'hFFFD;
        rom[81][23] = 16'h0009;
        rom[81][24] = 16'hFFF4;
        rom[81][25] = 16'h0000;
        rom[81][26] = 16'h0007;
        rom[81][27] = 16'h0008;
        rom[81][28] = 16'hFFE9;
        rom[81][29] = 16'hFFEB;
        rom[81][30] = 16'h0018;
        rom[81][31] = 16'hFFFE;
        rom[81][32] = 16'h0005;
        rom[81][33] = 16'h0006;
        rom[81][34] = 16'hFFC2;
        rom[81][35] = 16'h0010;
        rom[81][36] = 16'hFFD4;
        rom[81][37] = 16'h001C;
        rom[81][38] = 16'hFFD0;
        rom[81][39] = 16'h0026;
        rom[81][40] = 16'h0002;
        rom[81][41] = 16'hFFE0;
        rom[81][42] = 16'hFFC7;
        rom[81][43] = 16'h0014;
        rom[81][44] = 16'h0003;
        rom[81][45] = 16'hFFF4;
        rom[81][46] = 16'hFFFC;
        rom[81][47] = 16'hFFDF;
        rom[81][48] = 16'hFFF9;
        rom[81][49] = 16'h000C;
        rom[81][50] = 16'hFFD3;
        rom[81][51] = 16'h0033;
        rom[81][52] = 16'h0007;
        rom[81][53] = 16'hFFEB;
        rom[81][54] = 16'hFFF9;
        rom[81][55] = 16'h0020;
        rom[81][56] = 16'hFFC8;
        rom[81][57] = 16'h000C;
        rom[81][58] = 16'hFFEE;
        rom[81][59] = 16'hFFF4;
        rom[81][60] = 16'h0015;
        rom[81][61] = 16'h000E;
        rom[81][62] = 16'hFFEA;
        rom[81][63] = 16'h0041;
        rom[81][64] = 16'h000D;
        rom[81][65] = 16'hFFCD;
        rom[81][66] = 16'hFFD6;
        rom[81][67] = 16'h0010;
        rom[81][68] = 16'hFFEC;
        rom[81][69] = 16'hFFDB;
        rom[81][70] = 16'hFFD8;
        rom[81][71] = 16'h0007;
        rom[81][72] = 16'hFFDF;
        rom[81][73] = 16'hFFF2;
        rom[81][74] = 16'hFFCC;
        rom[81][75] = 16'hFFC8;
        rom[81][76] = 16'hFFC8;
        rom[81][77] = 16'hFFFC;
        rom[81][78] = 16'hFFF4;
        rom[81][79] = 16'hFFD5;
        rom[81][80] = 16'hFFE1;
        rom[81][81] = 16'h000B;
        rom[81][82] = 16'hFFEC;
        rom[81][83] = 16'h0003;
        rom[81][84] = 16'hFFCB;
        rom[81][85] = 16'hFFF2;
        rom[81][86] = 16'hFFF2;
        rom[81][87] = 16'h0006;
        rom[81][88] = 16'h0016;
        rom[81][89] = 16'hFFFE;
        rom[81][90] = 16'hFFE5;
        rom[81][91] = 16'hFFEA;
        rom[81][92] = 16'hFFF4;
        rom[81][93] = 16'h000A;
        rom[81][94] = 16'hFFDD;
        rom[81][95] = 16'h001B;
        rom[81][96] = 16'h001F;
        rom[81][97] = 16'h0016;
        rom[81][98] = 16'hFFE8;
        rom[81][99] = 16'h000C;
        rom[81][100] = 16'hFFF6;
        rom[81][101] = 16'h0016;
        rom[81][102] = 16'h0025;
        rom[81][103] = 16'h002A;
        rom[81][104] = 16'h0019;
        rom[81][105] = 16'h0036;
        rom[81][106] = 16'hFFDF;
        rom[81][107] = 16'hFFE3;
        rom[81][108] = 16'hFFF5;
        rom[81][109] = 16'hFFFC;
        rom[81][110] = 16'hFFE1;
        rom[81][111] = 16'hFFCD;
        rom[81][112] = 16'h0007;
        rom[81][113] = 16'h001D;
        rom[81][114] = 16'hFFFA;
        rom[81][115] = 16'hFFD0;
        rom[81][116] = 16'h000B;
        rom[81][117] = 16'hFFEA;
        rom[81][118] = 16'hFFF2;
        rom[81][119] = 16'hFFE3;
        rom[81][120] = 16'hFFFD;
        rom[81][121] = 16'hFFE0;
        rom[81][122] = 16'h0002;
        rom[81][123] = 16'hFFDD;
        rom[81][124] = 16'hFFE9;
        rom[81][125] = 16'h0012;
        rom[81][126] = 16'h000C;
        rom[81][127] = 16'hFFF4;
        rom[82][0] = 16'hFFDD;
        rom[82][1] = 16'hFFFF;
        rom[82][2] = 16'hFFFE;
        rom[82][3] = 16'hFFE8;
        rom[82][4] = 16'hFFEB;
        rom[82][5] = 16'hFFE4;
        rom[82][6] = 16'hFFEF;
        rom[82][7] = 16'hFFF4;
        rom[82][8] = 16'hFFB1;
        rom[82][9] = 16'hFFAB;
        rom[82][10] = 16'hFFEF;
        rom[82][11] = 16'h003D;
        rom[82][12] = 16'h0020;
        rom[82][13] = 16'hFFDD;
        rom[82][14] = 16'hFFC4;
        rom[82][15] = 16'h000A;
        rom[82][16] = 16'h0012;
        rom[82][17] = 16'hFFCD;
        rom[82][18] = 16'h002E;
        rom[82][19] = 16'h0001;
        rom[82][20] = 16'h0019;
        rom[82][21] = 16'hFFE3;
        rom[82][22] = 16'hFFD5;
        rom[82][23] = 16'hFFF6;
        rom[82][24] = 16'hFFF1;
        rom[82][25] = 16'hFFD7;
        rom[82][26] = 16'hFFFC;
        rom[82][27] = 16'hFFC3;
        rom[82][28] = 16'h001B;
        rom[82][29] = 16'hFFDD;
        rom[82][30] = 16'hFFF6;
        rom[82][31] = 16'hFFD6;
        rom[82][32] = 16'h0029;
        rom[82][33] = 16'hFFB5;
        rom[82][34] = 16'hFFDC;
        rom[82][35] = 16'h0000;
        rom[82][36] = 16'h0019;
        rom[82][37] = 16'hFFC8;
        rom[82][38] = 16'hFFBA;
        rom[82][39] = 16'hFFF2;
        rom[82][40] = 16'hFFD3;
        rom[82][41] = 16'h0024;
        rom[82][42] = 16'hFFCD;
        rom[82][43] = 16'h001B;
        rom[82][44] = 16'hFFF2;
        rom[82][45] = 16'h0019;
        rom[82][46] = 16'h002B;
        rom[82][47] = 16'hFFF2;
        rom[82][48] = 16'h0021;
        rom[82][49] = 16'h0006;
        rom[82][50] = 16'h0000;
        rom[82][51] = 16'hFFC9;
        rom[82][52] = 16'hFFEC;
        rom[82][53] = 16'hFFD6;
        rom[82][54] = 16'h0010;
        rom[82][55] = 16'hFFE1;
        rom[82][56] = 16'h000F;
        rom[82][57] = 16'hFFE6;
        rom[82][58] = 16'hFFF4;
        rom[82][59] = 16'h0004;
        rom[82][60] = 16'h0016;
        rom[82][61] = 16'h0001;
        rom[82][62] = 16'h001B;
        rom[82][63] = 16'h000B;
        rom[82][64] = 16'h0017;
        rom[82][65] = 16'h0016;
        rom[82][66] = 16'hFFC3;
        rom[82][67] = 16'hFFC4;
        rom[82][68] = 16'hFFE6;
        rom[82][69] = 16'hFFF7;
        rom[82][70] = 16'hFFC3;
        rom[82][71] = 16'hFFF7;
        rom[82][72] = 16'h0007;
        rom[82][73] = 16'hFFEA;
        rom[82][74] = 16'hFFF0;
        rom[82][75] = 16'hFFC0;
        rom[82][76] = 16'hFFF0;
        rom[82][77] = 16'hFFDE;
        rom[82][78] = 16'h0008;
        rom[82][79] = 16'hFFE1;
        rom[82][80] = 16'hFFE7;
        rom[82][81] = 16'h0033;
        rom[82][82] = 16'h0007;
        rom[82][83] = 16'hFFF3;
        rom[82][84] = 16'h0029;
        rom[82][85] = 16'hFFF0;
        rom[82][86] = 16'h0004;
        rom[82][87] = 16'hFFDC;
        rom[82][88] = 16'hFFDA;
        rom[82][89] = 16'h0018;
        rom[82][90] = 16'h0018;
        rom[82][91] = 16'hFFF4;
        rom[82][92] = 16'hFFE5;
        rom[82][93] = 16'h0015;
        rom[82][94] = 16'hFFE6;
        rom[82][95] = 16'h000E;
        rom[82][96] = 16'h0016;
        rom[82][97] = 16'h001C;
        rom[82][98] = 16'h000A;
        rom[82][99] = 16'h001B;
        rom[82][100] = 16'h000C;
        rom[82][101] = 16'h0021;
        rom[82][102] = 16'h0029;
        rom[82][103] = 16'hFFD8;
        rom[82][104] = 16'hFFC7;
        rom[82][105] = 16'hFFCB;
        rom[82][106] = 16'hFFD7;
        rom[82][107] = 16'h000E;
        rom[82][108] = 16'h0039;
        rom[82][109] = 16'h0013;
        rom[82][110] = 16'hFFFB;
        rom[82][111] = 16'h000B;
        rom[82][112] = 16'h000F;
        rom[82][113] = 16'hFFD4;
        rom[82][114] = 16'h0015;
        rom[82][115] = 16'h001F;
        rom[82][116] = 16'hFFEF;
        rom[82][117] = 16'h001F;
        rom[82][118] = 16'h0000;
        rom[82][119] = 16'h001D;
        rom[82][120] = 16'h0015;
        rom[82][121] = 16'hFFC1;
        rom[82][122] = 16'h000B;
        rom[82][123] = 16'hFFE7;
        rom[82][124] = 16'h0006;
        rom[82][125] = 16'hFFEC;
        rom[82][126] = 16'hFFEA;
        rom[82][127] = 16'hFFEF;
        rom[83][0] = 16'h0012;
        rom[83][1] = 16'h0019;
        rom[83][2] = 16'hFFC8;
        rom[83][3] = 16'hFFFB;
        rom[83][4] = 16'h0035;
        rom[83][5] = 16'hFFEA;
        rom[83][6] = 16'hFFE2;
        rom[83][7] = 16'h001C;
        rom[83][8] = 16'h002E;
        rom[83][9] = 16'h0000;
        rom[83][10] = 16'h0014;
        rom[83][11] = 16'h0021;
        rom[83][12] = 16'hFFF1;
        rom[83][13] = 16'h003C;
        rom[83][14] = 16'hFFE1;
        rom[83][15] = 16'hFFF6;
        rom[83][16] = 16'h000D;
        rom[83][17] = 16'hFFF7;
        rom[83][18] = 16'h001A;
        rom[83][19] = 16'hFFE9;
        rom[83][20] = 16'h0024;
        rom[83][21] = 16'h001E;
        rom[83][22] = 16'hFFD0;
        rom[83][23] = 16'hFFE1;
        rom[83][24] = 16'hFFEF;
        rom[83][25] = 16'hFFDE;
        rom[83][26] = 16'h0008;
        rom[83][27] = 16'hFFD0;
        rom[83][28] = 16'hFFEF;
        rom[83][29] = 16'h0011;
        rom[83][30] = 16'h002D;
        rom[83][31] = 16'h000C;
        rom[83][32] = 16'h0024;
        rom[83][33] = 16'h001D;
        rom[83][34] = 16'h0014;
        rom[83][35] = 16'h0015;
        rom[83][36] = 16'h002F;
        rom[83][37] = 16'h000F;
        rom[83][38] = 16'hFFD2;
        rom[83][39] = 16'hFFDE;
        rom[83][40] = 16'h000F;
        rom[83][41] = 16'hFFF4;
        rom[83][42] = 16'hFFF4;
        rom[83][43] = 16'hFFDC;
        rom[83][44] = 16'hFFC6;
        rom[83][45] = 16'hFFD0;
        rom[83][46] = 16'hFFF9;
        rom[83][47] = 16'hFFC4;
        rom[83][48] = 16'hFFC0;
        rom[83][49] = 16'hFFF9;
        rom[83][50] = 16'hFFC3;
        rom[83][51] = 16'hFFD7;
        rom[83][52] = 16'hFFC5;
        rom[83][53] = 16'hFFEB;
        rom[83][54] = 16'hFFFC;
        rom[83][55] = 16'hFFF0;
        rom[83][56] = 16'h001D;
        rom[83][57] = 16'hFFEC;
        rom[83][58] = 16'hFFD2;
        rom[83][59] = 16'h0023;
        rom[83][60] = 16'h0034;
        rom[83][61] = 16'hFFF7;
        rom[83][62] = 16'hFFE4;
        rom[83][63] = 16'hFFCB;
        rom[83][64] = 16'hFFFE;
        rom[83][65] = 16'h0038;
        rom[83][66] = 16'h000C;
        rom[83][67] = 16'h003F;
        rom[83][68] = 16'hFFE9;
        rom[83][69] = 16'hFFFE;
        rom[83][70] = 16'hFFF5;
        rom[83][71] = 16'hFFC5;
        rom[83][72] = 16'h001B;
        rom[83][73] = 16'hFFF5;
        rom[83][74] = 16'hFFF6;
        rom[83][75] = 16'h0007;
        rom[83][76] = 16'hFFE2;
        rom[83][77] = 16'h0011;
        rom[83][78] = 16'hFFB2;
        rom[83][79] = 16'hFFEF;
        rom[83][80] = 16'hFFD9;
        rom[83][81] = 16'h000B;
        rom[83][82] = 16'h0010;
        rom[83][83] = 16'h0001;
        rom[83][84] = 16'hFFF1;
        rom[83][85] = 16'h0000;
        rom[83][86] = 16'h0007;
        rom[83][87] = 16'hFFFD;
        rom[83][88] = 16'hFFBB;
        rom[83][89] = 16'hFFFD;
        rom[83][90] = 16'hFFFB;
        rom[83][91] = 16'hFFF9;
        rom[83][92] = 16'h000D;
        rom[83][93] = 16'hFFFF;
        rom[83][94] = 16'h0000;
        rom[83][95] = 16'hFFD6;
        rom[83][96] = 16'hFFDE;
        rom[83][97] = 16'hFFF7;
        rom[83][98] = 16'hFFE9;
        rom[83][99] = 16'h002D;
        rom[83][100] = 16'hFFC3;
        rom[83][101] = 16'hFFEF;
        rom[83][102] = 16'hFFEA;
        rom[83][103] = 16'h0002;
        rom[83][104] = 16'hFFDC;
        rom[83][105] = 16'hFFD7;
        rom[83][106] = 16'hFFD9;
        rom[83][107] = 16'hFFDE;
        rom[83][108] = 16'hFFFF;
        rom[83][109] = 16'hFFF6;
        rom[83][110] = 16'h0019;
        rom[83][111] = 16'hFFFC;
        rom[83][112] = 16'hFFCA;
        rom[83][113] = 16'hFFC3;
        rom[83][114] = 16'h0022;
        rom[83][115] = 16'h0028;
        rom[83][116] = 16'h0020;
        rom[83][117] = 16'h0006;
        rom[83][118] = 16'hFFE5;
        rom[83][119] = 16'hFFE7;
        rom[83][120] = 16'h002B;
        rom[83][121] = 16'hFFD5;
        rom[83][122] = 16'h000D;
        rom[83][123] = 16'h0016;
        rom[83][124] = 16'hFFE1;
        rom[83][125] = 16'hFFF0;
        rom[83][126] = 16'hFFBA;
        rom[83][127] = 16'hFFE2;
        rom[84][0] = 16'hFFF4;
        rom[84][1] = 16'hFFD4;
        rom[84][2] = 16'h0026;
        rom[84][3] = 16'hFFEB;
        rom[84][4] = 16'h001C;
        rom[84][5] = 16'h0002;
        rom[84][6] = 16'h0002;
        rom[84][7] = 16'hFFFD;
        rom[84][8] = 16'h0016;
        rom[84][9] = 16'h001F;
        rom[84][10] = 16'hFFF4;
        rom[84][11] = 16'hFFD8;
        rom[84][12] = 16'h000F;
        rom[84][13] = 16'hFFFE;
        rom[84][14] = 16'hFFEE;
        rom[84][15] = 16'hFFBD;
        rom[84][16] = 16'hFFF0;
        rom[84][17] = 16'h0000;
        rom[84][18] = 16'h0018;
        rom[84][19] = 16'hFFC4;
        rom[84][20] = 16'h0041;
        rom[84][21] = 16'hFFF9;
        rom[84][22] = 16'hFFF6;
        rom[84][23] = 16'hFFC4;
        rom[84][24] = 16'hFFEF;
        rom[84][25] = 16'h0015;
        rom[84][26] = 16'hFFC1;
        rom[84][27] = 16'h0011;
        rom[84][28] = 16'hFFF4;
        rom[84][29] = 16'h000C;
        rom[84][30] = 16'hFFD9;
        rom[84][31] = 16'h000E;
        rom[84][32] = 16'h000C;
        rom[84][33] = 16'hFFEA;
        rom[84][34] = 16'h0038;
        rom[84][35] = 16'h0029;
        rom[84][36] = 16'h000B;
        rom[84][37] = 16'hFFEF;
        rom[84][38] = 16'h0007;
        rom[84][39] = 16'h001E;
        rom[84][40] = 16'h001B;
        rom[84][41] = 16'hFFEE;
        rom[84][42] = 16'hFFEF;
        rom[84][43] = 16'hFFF6;
        rom[84][44] = 16'h0026;
        rom[84][45] = 16'h0014;
        rom[84][46] = 16'hFFE1;
        rom[84][47] = 16'hFFE8;
        rom[84][48] = 16'h0032;
        rom[84][49] = 16'hFFF4;
        rom[84][50] = 16'h0010;
        rom[84][51] = 16'h0012;
        rom[84][52] = 16'hFFE5;
        rom[84][53] = 16'hFFF2;
        rom[84][54] = 16'hFFF9;
        rom[84][55] = 16'h0015;
        rom[84][56] = 16'h001E;
        rom[84][57] = 16'h001B;
        rom[84][58] = 16'h000B;
        rom[84][59] = 16'h0024;
        rom[84][60] = 16'hFFEF;
        rom[84][61] = 16'hFFFB;
        rom[84][62] = 16'h0004;
        rom[84][63] = 16'h0022;
        rom[84][64] = 16'hFFF6;
        rom[84][65] = 16'hFFF5;
        rom[84][66] = 16'hFFFF;
        rom[84][67] = 16'hFFE4;
        rom[84][68] = 16'h0015;
        rom[84][69] = 16'hFFD2;
        rom[84][70] = 16'hFFE1;
        rom[84][71] = 16'hFFFA;
        rom[84][72] = 16'hFFF3;
        rom[84][73] = 16'h001C;
        rom[84][74] = 16'h000F;
        rom[84][75] = 16'h0007;
        rom[84][76] = 16'hFFFE;
        rom[84][77] = 16'h0019;
        rom[84][78] = 16'h0000;
        rom[84][79] = 16'hFFFC;
        rom[84][80] = 16'hFFD3;
        rom[84][81] = 16'hFFFE;
        rom[84][82] = 16'hFFFF;
        rom[84][83] = 16'h0016;
        rom[84][84] = 16'h000C;
        rom[84][85] = 16'hFFF9;
        rom[84][86] = 16'hFFF4;
        rom[84][87] = 16'h0002;
        rom[84][88] = 16'h000A;
        rom[84][89] = 16'h001C;
        rom[84][90] = 16'hFFFD;
        rom[84][91] = 16'hFFD9;
        rom[84][92] = 16'h0028;
        rom[84][93] = 16'h0002;
        rom[84][94] = 16'hFFEB;
        rom[84][95] = 16'h0007;
        rom[84][96] = 16'hFFF2;
        rom[84][97] = 16'h0008;
        rom[84][98] = 16'hFFB6;
        rom[84][99] = 16'hFFF4;
        rom[84][100] = 16'hFFED;
        rom[84][101] = 16'hFFE7;
        rom[84][102] = 16'h0024;
        rom[84][103] = 16'h0001;
        rom[84][104] = 16'hFFFE;
        rom[84][105] = 16'h0013;
        rom[84][106] = 16'h0008;
        rom[84][107] = 16'h0012;
        rom[84][108] = 16'hFFE5;
        rom[84][109] = 16'h0023;
        rom[84][110] = 16'hFFF7;
        rom[84][111] = 16'hFFD2;
        rom[84][112] = 16'hFFEB;
        rom[84][113] = 16'hFFF9;
        rom[84][114] = 16'hFFF9;
        rom[84][115] = 16'h001A;
        rom[84][116] = 16'hFFF0;
        rom[84][117] = 16'h000F;
        rom[84][118] = 16'hFFFA;
        rom[84][119] = 16'h0011;
        rom[84][120] = 16'hFFE5;
        rom[84][121] = 16'hFFC3;
        rom[84][122] = 16'hFFDB;
        rom[84][123] = 16'h0024;
        rom[84][124] = 16'h0009;
        rom[84][125] = 16'hFFFB;
        rom[84][126] = 16'hFFE9;
        rom[84][127] = 16'h0011;
        rom[85][0] = 16'hFFEF;
        rom[85][1] = 16'hFFFB;
        rom[85][2] = 16'hFFD7;
        rom[85][3] = 16'h0001;
        rom[85][4] = 16'h0002;
        rom[85][5] = 16'hFFFE;
        rom[85][6] = 16'h0030;
        rom[85][7] = 16'hFFB5;
        rom[85][8] = 16'h0034;
        rom[85][9] = 16'hFFCB;
        rom[85][10] = 16'h000A;
        rom[85][11] = 16'h0004;
        rom[85][12] = 16'hFFE8;
        rom[85][13] = 16'hFFED;
        rom[85][14] = 16'hFFE9;
        rom[85][15] = 16'h0005;
        rom[85][16] = 16'hFFFB;
        rom[85][17] = 16'hFFB5;
        rom[85][18] = 16'hFFF6;
        rom[85][19] = 16'h0017;
        rom[85][20] = 16'hFFF3;
        rom[85][21] = 16'hFFF9;
        rom[85][22] = 16'h0009;
        rom[85][23] = 16'h0016;
        rom[85][24] = 16'hFFC6;
        rom[85][25] = 16'h0028;
        rom[85][26] = 16'hFFE0;
        rom[85][27] = 16'hFFF7;
        rom[85][28] = 16'hFFF5;
        rom[85][29] = 16'hFFCE;
        rom[85][30] = 16'hFFC3;
        rom[85][31] = 16'h000D;
        rom[85][32] = 16'hFFE5;
        rom[85][33] = 16'hFFD5;
        rom[85][34] = 16'h0027;
        rom[85][35] = 16'hFFF4;
        rom[85][36] = 16'hFFF5;
        rom[85][37] = 16'hFFCF;
        rom[85][38] = 16'hFFD0;
        rom[85][39] = 16'hFFF3;
        rom[85][40] = 16'h0002;
        rom[85][41] = 16'h0015;
        rom[85][42] = 16'h000F;
        rom[85][43] = 16'hFFD5;
        rom[85][44] = 16'hFFF5;
        rom[85][45] = 16'h0024;
        rom[85][46] = 16'h0008;
        rom[85][47] = 16'h000B;
        rom[85][48] = 16'hFFE3;
        rom[85][49] = 16'h0004;
        rom[85][50] = 16'hFFEA;
        rom[85][51] = 16'hFFF4;
        rom[85][52] = 16'hFFFE;
        rom[85][53] = 16'h000B;
        rom[85][54] = 16'h002F;
        rom[85][55] = 16'hFFEF;
        rom[85][56] = 16'h000D;
        rom[85][57] = 16'h0014;
        rom[85][58] = 16'hFFEA;
        rom[85][59] = 16'h0016;
        rom[85][60] = 16'hFFE4;
        rom[85][61] = 16'hFFD8;
        rom[85][62] = 16'h002E;
        rom[85][63] = 16'h000F;
        rom[85][64] = 16'hFFA3;
        rom[85][65] = 16'hFFD3;
        rom[85][66] = 16'h001F;
        rom[85][67] = 16'h000C;
        rom[85][68] = 16'h001B;
        rom[85][69] = 16'h000F;
        rom[85][70] = 16'hFFE1;
        rom[85][71] = 16'h001E;
        rom[85][72] = 16'hFFCA;
        rom[85][73] = 16'h0007;
        rom[85][74] = 16'hFFF8;
        rom[85][75] = 16'hFFEF;
        rom[85][76] = 16'hFFD7;
        rom[85][77] = 16'hFFE0;
        rom[85][78] = 16'h0010;
        rom[85][79] = 16'hFFEA;
        rom[85][80] = 16'h001A;
        rom[85][81] = 16'h0016;
        rom[85][82] = 16'h000F;
        rom[85][83] = 16'h0016;
        rom[85][84] = 16'h0001;
        rom[85][85] = 16'hFFDE;
        rom[85][86] = 16'hFFEC;
        rom[85][87] = 16'hFFFF;
        rom[85][88] = 16'h0023;
        rom[85][89] = 16'h0023;
        rom[85][90] = 16'h0010;
        rom[85][91] = 16'h001F;
        rom[85][92] = 16'hFFEE;
        rom[85][93] = 16'h0000;
        rom[85][94] = 16'hFFF7;
        rom[85][95] = 16'hFFEF;
        rom[85][96] = 16'h000F;
        rom[85][97] = 16'h000B;
        rom[85][98] = 16'h0002;
        rom[85][99] = 16'h001B;
        rom[85][100] = 16'h001F;
        rom[85][101] = 16'h0005;
        rom[85][102] = 16'hFFF8;
        rom[85][103] = 16'h001D;
        rom[85][104] = 16'h0012;
        rom[85][105] = 16'h001C;
        rom[85][106] = 16'hFFEB;
        rom[85][107] = 16'h0023;
        rom[85][108] = 16'h0024;
        rom[85][109] = 16'hFFE3;
        rom[85][110] = 16'hFFFF;
        rom[85][111] = 16'h0015;
        rom[85][112] = 16'h0011;
        rom[85][113] = 16'h0007;
        rom[85][114] = 16'h0011;
        rom[85][115] = 16'hFFEC;
        rom[85][116] = 16'h0011;
        rom[85][117] = 16'h0009;
        rom[85][118] = 16'h002E;
        rom[85][119] = 16'h0002;
        rom[85][120] = 16'hFFC2;
        rom[85][121] = 16'h001B;
        rom[85][122] = 16'h0003;
        rom[85][123] = 16'hFFBA;
        rom[85][124] = 16'h002A;
        rom[85][125] = 16'h0001;
        rom[85][126] = 16'hFFD3;
        rom[85][127] = 16'h001F;
        rom[86][0] = 16'h0007;
        rom[86][1] = 16'hFFC8;
        rom[86][2] = 16'hFFD2;
        rom[86][3] = 16'h0027;
        rom[86][4] = 16'hFFE1;
        rom[86][5] = 16'hFFFB;
        rom[86][6] = 16'hFFE1;
        rom[86][7] = 16'h000D;
        rom[86][8] = 16'hFFDA;
        rom[86][9] = 16'h0030;
        rom[86][10] = 16'hFFEF;
        rom[86][11] = 16'hFFE0;
        rom[86][12] = 16'h0015;
        rom[86][13] = 16'h0007;
        rom[86][14] = 16'hFFEF;
        rom[86][15] = 16'h0019;
        rom[86][16] = 16'hFFF4;
        rom[86][17] = 16'hFFF2;
        rom[86][18] = 16'hFFDE;
        rom[86][19] = 16'hFFD2;
        rom[86][20] = 16'hFFE5;
        rom[86][21] = 16'hFFE5;
        rom[86][22] = 16'h0005;
        rom[86][23] = 16'hFFF9;
        rom[86][24] = 16'h000E;
        rom[86][25] = 16'hFFF6;
        rom[86][26] = 16'hFFB5;
        rom[86][27] = 16'h001B;
        rom[86][28] = 16'h0016;
        rom[86][29] = 16'h0011;
        rom[86][30] = 16'hFFE2;
        rom[86][31] = 16'h0002;
        rom[86][32] = 16'hFFB4;
        rom[86][33] = 16'h0000;
        rom[86][34] = 16'hFFDC;
        rom[86][35] = 16'h001F;
        rom[86][36] = 16'hFFD2;
        rom[86][37] = 16'hFFF8;
        rom[86][38] = 16'hFFCA;
        rom[86][39] = 16'h0010;
        rom[86][40] = 16'h002C;
        rom[86][41] = 16'hFFF9;
        rom[86][42] = 16'h002D;
        rom[86][43] = 16'hFFDC;
        rom[86][44] = 16'hFFD7;
        rom[86][45] = 16'h000D;
        rom[86][46] = 16'hFFEF;
        rom[86][47] = 16'h0033;
        rom[86][48] = 16'h0028;
        rom[86][49] = 16'hFFCB;
        rom[86][50] = 16'hFFD4;
        rom[86][51] = 16'hFFE8;
        rom[86][52] = 16'hFFB4;
        rom[86][53] = 16'h001D;
        rom[86][54] = 16'hFFFC;
        rom[86][55] = 16'hFFFE;
        rom[86][56] = 16'h0036;
        rom[86][57] = 16'hFFD2;
        rom[86][58] = 16'hFFFE;
        rom[86][59] = 16'hFFED;
        rom[86][60] = 16'hFFEA;
        rom[86][61] = 16'hFFF4;
        rom[86][62] = 16'h0029;
        rom[86][63] = 16'hFFF3;
        rom[86][64] = 16'h0005;
        rom[86][65] = 16'hFFF6;
        rom[86][66] = 16'hFFE5;
        rom[86][67] = 16'h0002;
        rom[86][68] = 16'h000B;
        rom[86][69] = 16'h0024;
        rom[86][70] = 16'hFFD2;
        rom[86][71] = 16'hFFD7;
        rom[86][72] = 16'hFFED;
        rom[86][73] = 16'hFFFC;
        rom[86][74] = 16'h0017;
        rom[86][75] = 16'h0017;
        rom[86][76] = 16'h0014;
        rom[86][77] = 16'h0008;
        rom[86][78] = 16'h0013;
        rom[86][79] = 16'h0003;
        rom[86][80] = 16'h0033;
        rom[86][81] = 16'hFFDF;
        rom[86][82] = 16'hFFBF;
        rom[86][83] = 16'hFFEF;
        rom[86][84] = 16'hFFE1;
        rom[86][85] = 16'h0028;
        rom[86][86] = 16'h001C;
        rom[86][87] = 16'h0007;
        rom[86][88] = 16'hFFAF;
        rom[86][89] = 16'hFFF9;
        rom[86][90] = 16'hFFC8;
        rom[86][91] = 16'hFFF3;
        rom[86][92] = 16'hFFFF;
        rom[86][93] = 16'h0014;
        rom[86][94] = 16'h0010;
        rom[86][95] = 16'h0016;
        rom[86][96] = 16'hFFFB;
        rom[86][97] = 16'hFFFA;
        rom[86][98] = 16'hFFE1;
        rom[86][99] = 16'hFFFB;
        rom[86][100] = 16'h0021;
        rom[86][101] = 16'h0008;
        rom[86][102] = 16'hFFD9;
        rom[86][103] = 16'h0004;
        rom[86][104] = 16'h0010;
        rom[86][105] = 16'hFFBA;
        rom[86][106] = 16'h001B;
        rom[86][107] = 16'h0018;
        rom[86][108] = 16'hFFCC;
        rom[86][109] = 16'h0023;
        rom[86][110] = 16'h0007;
        rom[86][111] = 16'hFFF3;
        rom[86][112] = 16'h0007;
        rom[86][113] = 16'hFFE4;
        rom[86][114] = 16'hFFFB;
        rom[86][115] = 16'hFFDF;
        rom[86][116] = 16'hFFF9;
        rom[86][117] = 16'h0001;
        rom[86][118] = 16'h0007;
        rom[86][119] = 16'hFFD0;
        rom[86][120] = 16'h0019;
        rom[86][121] = 16'h0024;
        rom[86][122] = 16'hFFEA;
        rom[86][123] = 16'hFFFC;
        rom[86][124] = 16'hFFD1;
        rom[86][125] = 16'h0022;
        rom[86][126] = 16'hFFDB;
        rom[86][127] = 16'hFFD7;
        rom[87][0] = 16'hFFEC;
        rom[87][1] = 16'h0005;
        rom[87][2] = 16'hFFE1;
        rom[87][3] = 16'hFFAC;
        rom[87][4] = 16'h0028;
        rom[87][5] = 16'hFFEE;
        rom[87][6] = 16'h0010;
        rom[87][7] = 16'h0016;
        rom[87][8] = 16'hFFA9;
        rom[87][9] = 16'hFFE1;
        rom[87][10] = 16'h0038;
        rom[87][11] = 16'hFFF1;
        rom[87][12] = 16'h0012;
        rom[87][13] = 16'hFFDF;
        rom[87][14] = 16'hFFFF;
        rom[87][15] = 16'hFFE0;
        rom[87][16] = 16'hFFF4;
        rom[87][17] = 16'h000E;
        rom[87][18] = 16'hFFCD;
        rom[87][19] = 16'h001F;
        rom[87][20] = 16'hFFB4;
        rom[87][21] = 16'h001A;
        rom[87][22] = 16'h0006;
        rom[87][23] = 16'hFFCD;
        rom[87][24] = 16'hFFEF;
        rom[87][25] = 16'hFFD2;
        rom[87][26] = 16'h0011;
        rom[87][27] = 16'h0013;
        rom[87][28] = 16'hFFE1;
        rom[87][29] = 16'h0020;
        rom[87][30] = 16'h0037;
        rom[87][31] = 16'hFFBE;
        rom[87][32] = 16'hFFDB;
        rom[87][33] = 16'h0008;
        rom[87][34] = 16'h0021;
        rom[87][35] = 16'hFFE8;
        rom[87][36] = 16'hFFE1;
        rom[87][37] = 16'h0001;
        rom[87][38] = 16'h0027;
        rom[87][39] = 16'h0002;
        rom[87][40] = 16'h0001;
        rom[87][41] = 16'h001F;
        rom[87][42] = 16'h002B;
        rom[87][43] = 16'hFFF2;
        rom[87][44] = 16'h0011;
        rom[87][45] = 16'hFFEB;
        rom[87][46] = 16'h0018;
        rom[87][47] = 16'hFFDC;
        rom[87][48] = 16'hFFF7;
        rom[87][49] = 16'hFFEF;
        rom[87][50] = 16'h001C;
        rom[87][51] = 16'h0024;
        rom[87][52] = 16'h001B;
        rom[87][53] = 16'hFFDC;
        rom[87][54] = 16'h0027;
        rom[87][55] = 16'h000C;
        rom[87][56] = 16'hFFED;
        rom[87][57] = 16'h0014;
        rom[87][58] = 16'h0022;
        rom[87][59] = 16'h000C;
        rom[87][60] = 16'h001A;
        rom[87][61] = 16'h0016;
        rom[87][62] = 16'hFFEA;
        rom[87][63] = 16'h0007;
        rom[87][64] = 16'hFFFC;
        rom[87][65] = 16'hFFDC;
        rom[87][66] = 16'hFFF9;
        rom[87][67] = 16'h0012;
        rom[87][68] = 16'hFFDF;
        rom[87][69] = 16'hFFCC;
        rom[87][70] = 16'hFFFD;
        rom[87][71] = 16'h0012;
        rom[87][72] = 16'h000F;
        rom[87][73] = 16'h0013;
        rom[87][74] = 16'h001B;
        rom[87][75] = 16'h0024;
        rom[87][76] = 16'h0016;
        rom[87][77] = 16'h003D;
        rom[87][78] = 16'h0000;
        rom[87][79] = 16'h002C;
        rom[87][80] = 16'hFFE9;
        rom[87][81] = 16'hFFF9;
        rom[87][82] = 16'h000F;
        rom[87][83] = 16'h0020;
        rom[87][84] = 16'hFFF8;
        rom[87][85] = 16'h001F;
        rom[87][86] = 16'hFFEB;
        rom[87][87] = 16'h0006;
        rom[87][88] = 16'hFFD2;
        rom[87][89] = 16'h001B;
        rom[87][90] = 16'hFFEB;
        rom[87][91] = 16'hFFFF;
        rom[87][92] = 16'h0000;
        rom[87][93] = 16'hFFB6;
        rom[87][94] = 16'h0008;
        rom[87][95] = 16'hFFD1;
        rom[87][96] = 16'hFFD7;
        rom[87][97] = 16'hFFEE;
        rom[87][98] = 16'hFFBA;
        rom[87][99] = 16'hFFFF;
        rom[87][100] = 16'hFFD0;
        rom[87][101] = 16'h002E;
        rom[87][102] = 16'h004A;
        rom[87][103] = 16'hFFFF;
        rom[87][104] = 16'hFFEF;
        rom[87][105] = 16'hFFDF;
        rom[87][106] = 16'h0004;
        rom[87][107] = 16'hFFE2;
        rom[87][108] = 16'hFFDC;
        rom[87][109] = 16'hFFA9;
        rom[87][110] = 16'hFFFE;
        rom[87][111] = 16'hFFD1;
        rom[87][112] = 16'h0021;
        rom[87][113] = 16'hFFE9;
        rom[87][114] = 16'hFFEF;
        rom[87][115] = 16'hFFED;
        rom[87][116] = 16'hFFF1;
        rom[87][117] = 16'hFFDC;
        rom[87][118] = 16'h0029;
        rom[87][119] = 16'h0005;
        rom[87][120] = 16'hFFFE;
        rom[87][121] = 16'hFFCB;
        rom[87][122] = 16'h000C;
        rom[87][123] = 16'hFFE2;
        rom[87][124] = 16'h0018;
        rom[87][125] = 16'h0033;
        rom[87][126] = 16'hFFF4;
        rom[87][127] = 16'h002A;
        rom[88][0] = 16'h001A;
        rom[88][1] = 16'h000D;
        rom[88][2] = 16'h002C;
        rom[88][3] = 16'hFFC3;
        rom[88][4] = 16'h0007;
        rom[88][5] = 16'hFFD4;
        rom[88][6] = 16'h001E;
        rom[88][7] = 16'h001C;
        rom[88][8] = 16'hFFD2;
        rom[88][9] = 16'hFFB3;
        rom[88][10] = 16'hFFAE;
        rom[88][11] = 16'h002F;
        rom[88][12] = 16'hFFE6;
        rom[88][13] = 16'h0010;
        rom[88][14] = 16'hFFD9;
        rom[88][15] = 16'h0000;
        rom[88][16] = 16'h0016;
        rom[88][17] = 16'h000A;
        rom[88][18] = 16'h0008;
        rom[88][19] = 16'hFFF9;
        rom[88][20] = 16'hFFFA;
        rom[88][21] = 16'h0049;
        rom[88][22] = 16'hFFF0;
        rom[88][23] = 16'hFFD4;
        rom[88][24] = 16'h000C;
        rom[88][25] = 16'h002B;
        rom[88][26] = 16'h0024;
        rom[88][27] = 16'hFFCD;
        rom[88][28] = 16'hFFBF;
        rom[88][29] = 16'h000C;
        rom[88][30] = 16'h0003;
        rom[88][31] = 16'h0029;
        rom[88][32] = 16'h000A;
        rom[88][33] = 16'hFFFE;
        rom[88][34] = 16'h0006;
        rom[88][35] = 16'hFFF3;
        rom[88][36] = 16'h0033;
        rom[88][37] = 16'hFFEE;
        rom[88][38] = 16'hFFBC;
        rom[88][39] = 16'hFFE1;
        rom[88][40] = 16'h0004;
        rom[88][41] = 16'hFFF9;
        rom[88][42] = 16'hFFF9;
        rom[88][43] = 16'hFFF4;
        rom[88][44] = 16'hFFF4;
        rom[88][45] = 16'hFFE1;
        rom[88][46] = 16'h0019;
        rom[88][47] = 16'hFFDC;
        rom[88][48] = 16'h0002;
        rom[88][49] = 16'hFFF9;
        rom[88][50] = 16'hFFF4;
        rom[88][51] = 16'h002A;
        rom[88][52] = 16'hFFFF;
        rom[88][53] = 16'hFFE3;
        rom[88][54] = 16'h001F;
        rom[88][55] = 16'hFFE0;
        rom[88][56] = 16'h001B;
        rom[88][57] = 16'hFFF5;
        rom[88][58] = 16'h000C;
        rom[88][59] = 16'hFFF9;
        rom[88][60] = 16'hFFF4;
        rom[88][61] = 16'h000D;
        rom[88][62] = 16'h000F;
        rom[88][63] = 16'hFFFE;
        rom[88][64] = 16'h0016;
        rom[88][65] = 16'h003A;
        rom[88][66] = 16'hFFF3;
        rom[88][67] = 16'hFFE2;
        rom[88][68] = 16'hFFFE;
        rom[88][69] = 16'hFFE9;
        rom[88][70] = 16'h0010;
        rom[88][71] = 16'h0024;
        rom[88][72] = 16'h003B;
        rom[88][73] = 16'hFFD8;
        rom[88][74] = 16'h0036;
        rom[88][75] = 16'hFFC6;
        rom[88][76] = 16'h000A;
        rom[88][77] = 16'hFFB2;
        rom[88][78] = 16'h0008;
        rom[88][79] = 16'h0034;
        rom[88][80] = 16'h0000;
        rom[88][81] = 16'h001E;
        rom[88][82] = 16'h0016;
        rom[88][83] = 16'hFFDF;
        rom[88][84] = 16'h0010;
        rom[88][85] = 16'hFFC6;
        rom[88][86] = 16'h0015;
        rom[88][87] = 16'hFFDA;
        rom[88][88] = 16'h0025;
        rom[88][89] = 16'h0005;
        rom[88][90] = 16'h0026;
        rom[88][91] = 16'h0018;
        rom[88][92] = 16'hFFE5;
        rom[88][93] = 16'hFFF2;
        rom[88][94] = 16'hFFFA;
        rom[88][95] = 16'hFFC5;
        rom[88][96] = 16'hFFF9;
        rom[88][97] = 16'h0031;
        rom[88][98] = 16'h002B;
        rom[88][99] = 16'hFFEE;
        rom[88][100] = 16'h000B;
        rom[88][101] = 16'h0011;
        rom[88][102] = 16'h001F;
        rom[88][103] = 16'hFFF8;
        rom[88][104] = 16'h0009;
        rom[88][105] = 16'hFFBD;
        rom[88][106] = 16'hFFF2;
        rom[88][107] = 16'h0012;
        rom[88][108] = 16'h003B;
        rom[88][109] = 16'hFFC8;
        rom[88][110] = 16'h001B;
        rom[88][111] = 16'h000C;
        rom[88][112] = 16'hFFDC;
        rom[88][113] = 16'hFFDE;
        rom[88][114] = 16'h001B;
        rom[88][115] = 16'h002F;
        rom[88][116] = 16'hFFEB;
        rom[88][117] = 16'hFFDE;
        rom[88][118] = 16'hFFF8;
        rom[88][119] = 16'hFFF2;
        rom[88][120] = 16'hFFF8;
        rom[88][121] = 16'hFFC3;
        rom[88][122] = 16'h0024;
        rom[88][123] = 16'hFFF3;
        rom[88][124] = 16'h000A;
        rom[88][125] = 16'h0001;
        rom[88][126] = 16'hFFD4;
        rom[88][127] = 16'hFFFF;
        rom[89][0] = 16'hFFE3;
        rom[89][1] = 16'h0010;
        rom[89][2] = 16'h0037;
        rom[89][3] = 16'h0000;
        rom[89][4] = 16'hFFD3;
        rom[89][5] = 16'hFFFF;
        rom[89][6] = 16'h0002;
        rom[89][7] = 16'hFFEA;
        rom[89][8] = 16'hFFF6;
        rom[89][9] = 16'hFFF1;
        rom[89][10] = 16'hFFE5;
        rom[89][11] = 16'h000F;
        rom[89][12] = 16'h0016;
        rom[89][13] = 16'hFFD3;
        rom[89][14] = 16'hFFED;
        rom[89][15] = 16'h002E;
        rom[89][16] = 16'hFFF9;
        rom[89][17] = 16'hFFA5;
        rom[89][18] = 16'hFFE1;
        rom[89][19] = 16'hFFF4;
        rom[89][20] = 16'hFFE1;
        rom[89][21] = 16'h0014;
        rom[89][22] = 16'hFFCD;
        rom[89][23] = 16'hFFEE;
        rom[89][24] = 16'h0031;
        rom[89][25] = 16'hFFD2;
        rom[89][26] = 16'hFFE8;
        rom[89][27] = 16'hFFE8;
        rom[89][28] = 16'h0024;
        rom[89][29] = 16'hFFF1;
        rom[89][30] = 16'hFFEC;
        rom[89][31] = 16'hFFDA;
        rom[89][32] = 16'hFFE6;
        rom[89][33] = 16'hFFEA;
        rom[89][34] = 16'hFFA4;
        rom[89][35] = 16'h0013;
        rom[89][36] = 16'hFFF6;
        rom[89][37] = 16'hFFF2;
        rom[89][38] = 16'hFFFC;
        rom[89][39] = 16'hFFF7;
        rom[89][40] = 16'hFFAA;
        rom[89][41] = 16'h0000;
        rom[89][42] = 16'hFFD2;
        rom[89][43] = 16'h001F;
        rom[89][44] = 16'hFFFA;
        rom[89][45] = 16'hFFEF;
        rom[89][46] = 16'h000C;
        rom[89][47] = 16'h0010;
        rom[89][48] = 16'hFFFD;
        rom[89][49] = 16'hFFF5;
        rom[89][50] = 16'h002F;
        rom[89][51] = 16'hFFD1;
        rom[89][52] = 16'hFFFA;
        rom[89][53] = 16'h000F;
        rom[89][54] = 16'h0011;
        rom[89][55] = 16'h0011;
        rom[89][56] = 16'h0011;
        rom[89][57] = 16'hFFD5;
        rom[89][58] = 16'h0011;
        rom[89][59] = 16'hFFEF;
        rom[89][60] = 16'hFFEF;
        rom[89][61] = 16'h001B;
        rom[89][62] = 16'h0023;
        rom[89][63] = 16'hFFEB;
        rom[89][64] = 16'hFFFB;
        rom[89][65] = 16'hFFF1;
        rom[89][66] = 16'h001F;
        rom[89][67] = 16'h0011;
        rom[89][68] = 16'hFFCA;
        rom[89][69] = 16'h0016;
        rom[89][70] = 16'h000C;
        rom[89][71] = 16'h0019;
        rom[89][72] = 16'h0007;
        rom[89][73] = 16'hFFEA;
        rom[89][74] = 16'hFFB2;
        rom[89][75] = 16'h0008;
        rom[89][76] = 16'hFFFC;
        rom[89][77] = 16'hFFBE;
        rom[89][78] = 16'hFFEB;
        rom[89][79] = 16'hFFE5;
        rom[89][80] = 16'hFFFD;
        rom[89][81] = 16'h001C;
        rom[89][82] = 16'hFFFA;
        rom[89][83] = 16'h0017;
        rom[89][84] = 16'h000C;
        rom[89][85] = 16'hFFEE;
        rom[89][86] = 16'h0003;
        rom[89][87] = 16'hFFE8;
        rom[89][88] = 16'hFFCA;
        rom[89][89] = 16'h0006;
        rom[89][90] = 16'h0002;
        rom[89][91] = 16'hFFF0;
        rom[89][92] = 16'hFFE5;
        rom[89][93] = 16'hFFFD;
        rom[89][94] = 16'hFFC4;
        rom[89][95] = 16'hFFCE;
        rom[89][96] = 16'hFFFB;
        rom[89][97] = 16'hFFEB;
        rom[89][98] = 16'h0011;
        rom[89][99] = 16'h0009;
        rom[89][100] = 16'hFFFE;
        rom[89][101] = 16'hFFD3;
        rom[89][102] = 16'hFFD0;
        rom[89][103] = 16'hFFD4;
        rom[89][104] = 16'hFFDC;
        rom[89][105] = 16'hFFCD;
        rom[89][106] = 16'hFFE7;
        rom[89][107] = 16'h001B;
        rom[89][108] = 16'hFFFA;
        rom[89][109] = 16'h0031;
        rom[89][110] = 16'h0008;
        rom[89][111] = 16'h0022;
        rom[89][112] = 16'hFFFE;
        rom[89][113] = 16'h001B;
        rom[89][114] = 16'hFFFB;
        rom[89][115] = 16'hFFF4;
        rom[89][116] = 16'h0004;
        rom[89][117] = 16'hFFD1;
        rom[89][118] = 16'hFFF7;
        rom[89][119] = 16'h0039;
        rom[89][120] = 16'hFFE8;
        rom[89][121] = 16'hFFFF;
        rom[89][122] = 16'hFFE4;
        rom[89][123] = 16'hFFF7;
        rom[89][124] = 16'h0017;
        rom[89][125] = 16'hFFF1;
        rom[89][126] = 16'hFFF4;
        rom[89][127] = 16'h0004;
        rom[90][0] = 16'h000B;
        rom[90][1] = 16'h001C;
        rom[90][2] = 16'hFFEE;
        rom[90][3] = 16'hFFF2;
        rom[90][4] = 16'hFFE6;
        rom[90][5] = 16'h0031;
        rom[90][6] = 16'hFFE5;
        rom[90][7] = 16'h000E;
        rom[90][8] = 16'hFFBE;
        rom[90][9] = 16'h0008;
        rom[90][10] = 16'h0007;
        rom[90][11] = 16'h0009;
        rom[90][12] = 16'hFFF3;
        rom[90][13] = 16'h0024;
        rom[90][14] = 16'hFFAB;
        rom[90][15] = 16'hFFFE;
        rom[90][16] = 16'h0002;
        rom[90][17] = 16'h004B;
        rom[90][18] = 16'hFFEC;
        rom[90][19] = 16'hFFE8;
        rom[90][20] = 16'hFFF8;
        rom[90][21] = 16'h001F;
        rom[90][22] = 16'h0002;
        rom[90][23] = 16'hFFF8;
        rom[90][24] = 16'hFFE8;
        rom[90][25] = 16'hFFF4;
        rom[90][26] = 16'h0006;
        rom[90][27] = 16'h000B;
        rom[90][28] = 16'hFFBC;
        rom[90][29] = 16'hFFEA;
        rom[90][30] = 16'h0012;
        rom[90][31] = 16'hFFE0;
        rom[90][32] = 16'h003F;
        rom[90][33] = 16'hFFF8;
        rom[90][34] = 16'hFFE2;
        rom[90][35] = 16'h000E;
        rom[90][36] = 16'h003B;
        rom[90][37] = 16'hFFE1;
        rom[90][38] = 16'h001D;
        rom[90][39] = 16'hFFE8;
        rom[90][40] = 16'hFFF7;
        rom[90][41] = 16'h0016;
        rom[90][42] = 16'h0029;
        rom[90][43] = 16'hFFCF;
        rom[90][44] = 16'h0008;
        rom[90][45] = 16'h0011;
        rom[90][46] = 16'hFFFE;
        rom[90][47] = 16'h0006;
        rom[90][48] = 16'h0020;
        rom[90][49] = 16'h0028;
        rom[90][50] = 16'hFFF7;
        rom[90][51] = 16'h002F;
        rom[90][52] = 16'hFFB5;
        rom[90][53] = 16'hFFE1;
        rom[90][54] = 16'hFFDD;
        rom[90][55] = 16'h000F;
        rom[90][56] = 16'h0024;
        rom[90][57] = 16'hFFE3;
        rom[90][58] = 16'hFFDF;
        rom[90][59] = 16'hFFEE;
        rom[90][60] = 16'hFFE5;
        rom[90][61] = 16'h0019;
        rom[90][62] = 16'hFFE8;
        rom[90][63] = 16'h0002;
        rom[90][64] = 16'h0016;
        rom[90][65] = 16'hFFEF;
        rom[90][66] = 16'hFFCF;
        rom[90][67] = 16'h0002;
        rom[90][68] = 16'hFFE1;
        rom[90][69] = 16'h0002;
        rom[90][70] = 16'h001A;
        rom[90][71] = 16'hFFE1;
        rom[90][72] = 16'h001A;
        rom[90][73] = 16'hFFF9;
        rom[90][74] = 16'hFFFC;
        rom[90][75] = 16'hFFE8;
        rom[90][76] = 16'hFFF5;
        rom[90][77] = 16'hFFFD;
        rom[90][78] = 16'h0005;
        rom[90][79] = 16'h0007;
        rom[90][80] = 16'hFFFB;
        rom[90][81] = 16'h0018;
        rom[90][82] = 16'h0027;
        rom[90][83] = 16'hFFF4;
        rom[90][84] = 16'h0021;
        rom[90][85] = 16'hFFFB;
        rom[90][86] = 16'h0010;
        rom[90][87] = 16'h0004;
        rom[90][88] = 16'h0001;
        rom[90][89] = 16'h0000;
        rom[90][90] = 16'h000F;
        rom[90][91] = 16'h0002;
        rom[90][92] = 16'hFFAB;
        rom[90][93] = 16'hFFD2;
        rom[90][94] = 16'hFFBE;
        rom[90][95] = 16'h0017;
        rom[90][96] = 16'hFFF9;
        rom[90][97] = 16'hFFCD;
        rom[90][98] = 16'hFFC6;
        rom[90][99] = 16'h001C;
        rom[90][100] = 16'hFFFB;
        rom[90][101] = 16'h0035;
        rom[90][102] = 16'hFFEA;
        rom[90][103] = 16'hFFD3;
        rom[90][104] = 16'h003D;
        rom[90][105] = 16'hFFEF;
        rom[90][106] = 16'hFFF4;
        rom[90][107] = 16'h0017;
        rom[90][108] = 16'h0002;
        rom[90][109] = 16'h0028;
        rom[90][110] = 16'h0008;
        rom[90][111] = 16'hFFE5;
        rom[90][112] = 16'h0010;
        rom[90][113] = 16'h0020;
        rom[90][114] = 16'hFFD0;
        rom[90][115] = 16'hFFF7;
        rom[90][116] = 16'hFFDD;
        rom[90][117] = 16'h0006;
        rom[90][118] = 16'h0024;
        rom[90][119] = 16'h0017;
        rom[90][120] = 16'hFFEC;
        rom[90][121] = 16'hFFCF;
        rom[90][122] = 16'hFFE6;
        rom[90][123] = 16'hFFFA;
        rom[90][124] = 16'hFFD9;
        rom[90][125] = 16'hFFF8;
        rom[90][126] = 16'hFFE0;
        rom[90][127] = 16'h000A;
        rom[91][0] = 16'h0012;
        rom[91][1] = 16'hFFD1;
        rom[91][2] = 16'h000F;
        rom[91][3] = 16'hFFFB;
        rom[91][4] = 16'hFFFE;
        rom[91][5] = 16'hFFFF;
        rom[91][6] = 16'h0018;
        rom[91][7] = 16'hFFB1;
        rom[91][8] = 16'h0009;
        rom[91][9] = 16'h0016;
        rom[91][10] = 16'h002C;
        rom[91][11] = 16'h0013;
        rom[91][12] = 16'h0018;
        rom[91][13] = 16'hFFC0;
        rom[91][14] = 16'h0021;
        rom[91][15] = 16'hFFD9;
        rom[91][16] = 16'h0016;
        rom[91][17] = 16'hFFDE;
        rom[91][18] = 16'h001E;
        rom[91][19] = 16'hFFE5;
        rom[91][20] = 16'hFFFE;
        rom[91][21] = 16'hFFE1;
        rom[91][22] = 16'hFFE9;
        rom[91][23] = 16'h0007;
        rom[91][24] = 16'hFFEF;
        rom[91][25] = 16'hFFF7;
        rom[91][26] = 16'h000B;
        rom[91][27] = 16'hFFF7;
        rom[91][28] = 16'hFFEE;
        rom[91][29] = 16'hFFC7;
        rom[91][30] = 16'h0016;
        rom[91][31] = 16'hFFEF;
        rom[91][32] = 16'hFFF6;
        rom[91][33] = 16'hFFA2;
        rom[91][34] = 16'hFFD0;
        rom[91][35] = 16'hFFC8;
        rom[91][36] = 16'hFFE5;
        rom[91][37] = 16'hFFCF;
        rom[91][38] = 16'hFFE5;
        rom[91][39] = 16'h0002;
        rom[91][40] = 16'hFFFE;
        rom[91][41] = 16'hFFFA;
        rom[91][42] = 16'h002C;
        rom[91][43] = 16'hFFF1;
        rom[91][44] = 16'h0038;
        rom[91][45] = 16'hFFE6;
        rom[91][46] = 16'hFFE2;
        rom[91][47] = 16'hFFF9;
        rom[91][48] = 16'hFFE3;
        rom[91][49] = 16'hFFD2;
        rom[91][50] = 16'h0002;
        rom[91][51] = 16'h0035;
        rom[91][52] = 16'hFFEB;
        rom[91][53] = 16'hFFF0;
        rom[91][54] = 16'h001D;
        rom[91][55] = 16'h0025;
        rom[91][56] = 16'hFFEF;
        rom[91][57] = 16'h0000;
        rom[91][58] = 16'h0015;
        rom[91][59] = 16'h001C;
        rom[91][60] = 16'h0016;
        rom[91][61] = 16'hFFBB;
        rom[91][62] = 16'hFFFF;
        rom[91][63] = 16'h0009;
        rom[91][64] = 16'hFFC7;
        rom[91][65] = 16'hFFBA;
        rom[91][66] = 16'h000A;
        rom[91][67] = 16'h000C;
        rom[91][68] = 16'hFFF4;
        rom[91][69] = 16'h000E;
        rom[91][70] = 16'hFFDA;
        rom[91][71] = 16'hFFEC;
        rom[91][72] = 16'h0002;
        rom[91][73] = 16'hFFEB;
        rom[91][74] = 16'h0016;
        rom[91][75] = 16'hFFE1;
        rom[91][76] = 16'hFFDC;
        rom[91][77] = 16'h0026;
        rom[91][78] = 16'h0029;
        rom[91][79] = 16'hFFE7;
        rom[91][80] = 16'h0018;
        rom[91][81] = 16'hFFCF;
        rom[91][82] = 16'hFFE0;
        rom[91][83] = 16'h0028;
        rom[91][84] = 16'hFFB4;
        rom[91][85] = 16'hFFFE;
        rom[91][86] = 16'h0016;
        rom[91][87] = 16'h0003;
        rom[91][88] = 16'h0007;
        rom[91][89] = 16'h000E;
        rom[91][90] = 16'hFFEE;
        rom[91][91] = 16'h0016;
        rom[91][92] = 16'h0009;
        rom[91][93] = 16'h0004;
        rom[91][94] = 16'hFFF4;
        rom[91][95] = 16'h0007;
        rom[91][96] = 16'hFFEE;
        rom[91][97] = 16'h0017;
        rom[91][98] = 16'h000E;
        rom[91][99] = 16'hFFC3;
        rom[91][100] = 16'hFFFF;
        rom[91][101] = 16'hFFE5;
        rom[91][102] = 16'hFFDE;
        rom[91][103] = 16'h0004;
        rom[91][104] = 16'h000B;
        rom[91][105] = 16'h0011;
        rom[91][106] = 16'h0000;
        rom[91][107] = 16'hFFFF;
        rom[91][108] = 16'hFFD9;
        rom[91][109] = 16'hFFE3;
        rom[91][110] = 16'hFFCF;
        rom[91][111] = 16'h0007;
        rom[91][112] = 16'hFFEA;
        rom[91][113] = 16'h001D;
        rom[91][114] = 16'hFFEC;
        rom[91][115] = 16'h0012;
        rom[91][116] = 16'hFFB2;
        rom[91][117] = 16'h0016;
        rom[91][118] = 16'h002A;
        rom[91][119] = 16'hFFE4;
        rom[91][120] = 16'hFFEA;
        rom[91][121] = 16'h0014;
        rom[91][122] = 16'h004B;
        rom[91][123] = 16'hFFE9;
        rom[91][124] = 16'h0011;
        rom[91][125] = 16'h0015;
        rom[91][126] = 16'hFFE5;
        rom[91][127] = 16'h000F;
        rom[92][0] = 16'hFFD7;
        rom[92][1] = 16'h0006;
        rom[92][2] = 16'h000C;
        rom[92][3] = 16'h002D;
        rom[92][4] = 16'hFFFF;
        rom[92][5] = 16'hFFED;
        rom[92][6] = 16'hFFCB;
        rom[92][7] = 16'hFFF8;
        rom[92][8] = 16'hFFEE;
        rom[92][9] = 16'h001B;
        rom[92][10] = 16'h0038;
        rom[92][11] = 16'h0006;
        rom[92][12] = 16'hFFF5;
        rom[92][13] = 16'hFFF8;
        rom[92][14] = 16'hFFF1;
        rom[92][15] = 16'hFFEA;
        rom[92][16] = 16'hFFEA;
        rom[92][17] = 16'h001F;
        rom[92][18] = 16'hFFF3;
        rom[92][19] = 16'h0007;
        rom[92][20] = 16'h0016;
        rom[92][21] = 16'hFFDD;
        rom[92][22] = 16'hFFF9;
        rom[92][23] = 16'h0013;
        rom[92][24] = 16'hFFEF;
        rom[92][25] = 16'hFFD0;
        rom[92][26] = 16'hFFF4;
        rom[92][27] = 16'h0016;
        rom[92][28] = 16'h002E;
        rom[92][29] = 16'h0000;
        rom[92][30] = 16'hFFFE;
        rom[92][31] = 16'hFFE0;
        rom[92][32] = 16'h0001;
        rom[92][33] = 16'hFFEF;
        rom[92][34] = 16'hFFFA;
        rom[92][35] = 16'h0001;
        rom[92][36] = 16'hFFD9;
        rom[92][37] = 16'h0009;
        rom[92][38] = 16'hFFEE;
        rom[92][39] = 16'hFFCF;
        rom[92][40] = 16'h0000;
        rom[92][41] = 16'hFFC3;
        rom[92][42] = 16'h0007;
        rom[92][43] = 16'h0010;
        rom[92][44] = 16'hFFF2;
        rom[92][45] = 16'h0024;
        rom[92][46] = 16'hFFEB;
        rom[92][47] = 16'hFFF7;
        rom[92][48] = 16'hFFF3;
        rom[92][49] = 16'hFFB4;
        rom[92][50] = 16'hFFFA;
        rom[92][51] = 16'h0000;
        rom[92][52] = 16'hFFF8;
        rom[92][53] = 16'h0016;
        rom[92][54] = 16'hFFF5;
        rom[92][55] = 16'hFFC8;
        rom[92][56] = 16'h0006;
        rom[92][57] = 16'hFFF8;
        rom[92][58] = 16'h0001;
        rom[92][59] = 16'h0027;
        rom[92][60] = 16'hFFE2;
        rom[92][61] = 16'h0018;
        rom[92][62] = 16'hFFE1;
        rom[92][63] = 16'hFFF9;
        rom[92][64] = 16'hFFA6;
        rom[92][65] = 16'hFFD5;
        rom[92][66] = 16'hFFEB;
        rom[92][67] = 16'h0003;
        rom[92][68] = 16'hFFBA;
        rom[92][69] = 16'hFFFF;
        rom[92][70] = 16'h0009;
        rom[92][71] = 16'h0010;
        rom[92][72] = 16'hFFF5;
        rom[92][73] = 16'hFFF1;
        rom[92][74] = 16'hFFE2;
        rom[92][75] = 16'hFFF8;
        rom[92][76] = 16'h0028;
        rom[92][77] = 16'h0005;
        rom[92][78] = 16'hFFCF;
        rom[92][79] = 16'h0018;
        rom[92][80] = 16'hFFE0;
        rom[92][81] = 16'hFFEE;
        rom[92][82] = 16'h0046;
        rom[92][83] = 16'hFFF6;
        rom[92][84] = 16'hFFF9;
        rom[92][85] = 16'hFFF4;
        rom[92][86] = 16'hFFF4;
        rom[92][87] = 16'h0010;
        rom[92][88] = 16'hFFCD;
        rom[92][89] = 16'hFFE1;
        rom[92][90] = 16'h0027;
        rom[92][91] = 16'h000C;
        rom[92][92] = 16'hFFF1;
        rom[92][93] = 16'hFFEA;
        rom[92][94] = 16'h001B;
        rom[92][95] = 16'h000F;
        rom[92][96] = 16'hFFE5;
        rom[92][97] = 16'hFFB8;
        rom[92][98] = 16'hFFE8;
        rom[92][99] = 16'hFFE4;
        rom[92][100] = 16'hFFED;
        rom[92][101] = 16'hFFBF;
        rom[92][102] = 16'hFFD7;
        rom[92][103] = 16'h0014;
        rom[92][104] = 16'h0024;
        rom[92][105] = 16'hFFF1;
        rom[92][106] = 16'h0028;
        rom[92][107] = 16'h002B;
        rom[92][108] = 16'hFFCD;
        rom[92][109] = 16'hFFF3;
        rom[92][110] = 16'h0021;
        rom[92][111] = 16'hFFEE;
        rom[92][112] = 16'h0006;
        rom[92][113] = 16'h0060;
        rom[92][114] = 16'h0018;
        rom[92][115] = 16'hFFE5;
        rom[92][116] = 16'h0010;
        rom[92][117] = 16'hFFDC;
        rom[92][118] = 16'h0004;
        rom[92][119] = 16'hFFEF;
        rom[92][120] = 16'h000C;
        rom[92][121] = 16'h0007;
        rom[92][122] = 16'h001A;
        rom[92][123] = 16'h0007;
        rom[92][124] = 16'hFFEA;
        rom[92][125] = 16'h0011;
        rom[92][126] = 16'h001A;
        rom[92][127] = 16'h0012;
        rom[93][0] = 16'hFFCE;
        rom[93][1] = 16'h0008;
        rom[93][2] = 16'h0002;
        rom[93][3] = 16'h0019;
        rom[93][4] = 16'hFFF4;
        rom[93][5] = 16'hFFF9;
        rom[93][6] = 16'h000C;
        rom[93][7] = 16'hFFFB;
        rom[93][8] = 16'h0019;
        rom[93][9] = 16'h0029;
        rom[93][10] = 16'hFFF2;
        rom[93][11] = 16'hFFF7;
        rom[93][12] = 16'h001D;
        rom[93][13] = 16'h0003;
        rom[93][14] = 16'hFFDE;
        rom[93][15] = 16'h002C;
        rom[93][16] = 16'hFFF2;
        rom[93][17] = 16'h0018;
        rom[93][18] = 16'hFFF1;
        rom[93][19] = 16'h002F;
        rom[93][20] = 16'hFFE3;
        rom[93][21] = 16'h000B;
        rom[93][22] = 16'hFFF8;
        rom[93][23] = 16'h0009;
        rom[93][24] = 16'h000C;
        rom[93][25] = 16'hFFF5;
        rom[93][26] = 16'hFFF8;
        rom[93][27] = 16'hFFEA;
        rom[93][28] = 16'h001E;
        rom[93][29] = 16'h000E;
        rom[93][30] = 16'hFFCB;
        rom[93][31] = 16'hFFB1;
        rom[93][32] = 16'hFFDB;
        rom[93][33] = 16'hFFE9;
        rom[93][34] = 16'h0005;
        rom[93][35] = 16'hFFEA;
        rom[93][36] = 16'hFFED;
        rom[93][37] = 16'h0009;
        rom[93][38] = 16'h004C;
        rom[93][39] = 16'h000E;
        rom[93][40] = 16'hFFFC;
        rom[93][41] = 16'h0009;
        rom[93][42] = 16'hFFE5;
        rom[93][43] = 16'hFFF4;
        rom[93][44] = 16'hFFEA;
        rom[93][45] = 16'hFFFB;
        rom[93][46] = 16'hFFE3;
        rom[93][47] = 16'hFFF4;
        rom[93][48] = 16'hFFE8;
        rom[93][49] = 16'hFFEC;
        rom[93][50] = 16'hFFE5;
        rom[93][51] = 16'hFFA3;
        rom[93][52] = 16'hFFFD;
        rom[93][53] = 16'hFFEA;
        rom[93][54] = 16'h0004;
        rom[93][55] = 16'h0000;
        rom[93][56] = 16'h000D;
        rom[93][57] = 16'hFFE9;
        rom[93][58] = 16'hFFFD;
        rom[93][59] = 16'hFFDC;
        rom[93][60] = 16'hFFDE;
        rom[93][61] = 16'h0029;
        rom[93][62] = 16'hFFF5;
        rom[93][63] = 16'h0000;
        rom[93][64] = 16'h001A;
        rom[93][65] = 16'hFFC9;
        rom[93][66] = 16'h0002;
        rom[93][67] = 16'h0007;
        rom[93][68] = 16'h0002;
        rom[93][69] = 16'h001F;
        rom[93][70] = 16'hFFDD;
        rom[93][71] = 16'hFFC9;
        rom[93][72] = 16'hFFC0;
        rom[93][73] = 16'h0013;
        rom[93][74] = 16'hFFCF;
        rom[93][75] = 16'h0002;
        rom[93][76] = 16'h0022;
        rom[93][77] = 16'hFFDC;
        rom[93][78] = 16'h000C;
        rom[93][79] = 16'hFFD6;
        rom[93][80] = 16'hFFFC;
        rom[93][81] = 16'h0027;
        rom[93][82] = 16'h000F;
        rom[93][83] = 16'h000B;
        rom[93][84] = 16'hFFEA;
        rom[93][85] = 16'h005F;
        rom[93][86] = 16'hFFF9;
        rom[93][87] = 16'hFFF9;
        rom[93][88] = 16'h0004;
        rom[93][89] = 16'hFFF4;
        rom[93][90] = 16'hFFEC;
        rom[93][91] = 16'hFFDB;
        rom[93][92] = 16'hFFDF;
        rom[93][93] = 16'h000F;
        rom[93][94] = 16'hFFF0;
        rom[93][95] = 16'hFFF4;
        rom[93][96] = 16'hFFFB;
        rom[93][97] = 16'h0027;
        rom[93][98] = 16'h000B;
        rom[93][99] = 16'h0023;
        rom[93][100] = 16'h0028;
        rom[93][101] = 16'hFFF6;
        rom[93][102] = 16'h0016;
        rom[93][103] = 16'hFFEE;
        rom[93][104] = 16'hFFB0;
        rom[93][105] = 16'h0013;
        rom[93][106] = 16'h0016;
        rom[93][107] = 16'hFFF8;
        rom[93][108] = 16'hFFEB;
        rom[93][109] = 16'hFFFC;
        rom[93][110] = 16'hFFFE;
        rom[93][111] = 16'hFFEC;
        rom[93][112] = 16'hFFE2;
        rom[93][113] = 16'h001B;
        rom[93][114] = 16'h000F;
        rom[93][115] = 16'hFFFC;
        rom[93][116] = 16'hFFE9;
        rom[93][117] = 16'hFFDA;
        rom[93][118] = 16'h0004;
        rom[93][119] = 16'h004D;
        rom[93][120] = 16'hFFE9;
        rom[93][121] = 16'h0006;
        rom[93][122] = 16'hFFE5;
        rom[93][123] = 16'hFFC6;
        rom[93][124] = 16'hFFFA;
        rom[93][125] = 16'hFFC4;
        rom[93][126] = 16'hFFE5;
        rom[93][127] = 16'hFFE1;
        rom[94][0] = 16'h000B;
        rom[94][1] = 16'hFFE0;
        rom[94][2] = 16'hFFF8;
        rom[94][3] = 16'h001A;
        rom[94][4] = 16'hFFE4;
        rom[94][5] = 16'hFFF3;
        rom[94][6] = 16'h001F;
        rom[94][7] = 16'hFFD7;
        rom[94][8] = 16'hFFF2;
        rom[94][9] = 16'hFFE8;
        rom[94][10] = 16'hFFE1;
        rom[94][11] = 16'hFFED;
        rom[94][12] = 16'hFFFC;
        rom[94][13] = 16'hFFF5;
        rom[94][14] = 16'hFFD8;
        rom[94][15] = 16'hFFE6;
        rom[94][16] = 16'hFFF1;
        rom[94][17] = 16'hFFD7;
        rom[94][18] = 16'hFFDB;
        rom[94][19] = 16'hFFE0;
        rom[94][20] = 16'hFFEA;
        rom[94][21] = 16'hFFF9;
        rom[94][22] = 16'h002E;
        rom[94][23] = 16'hFFF6;
        rom[94][24] = 16'hFFF4;
        rom[94][25] = 16'h0015;
        rom[94][26] = 16'hFFB5;
        rom[94][27] = 16'h001B;
        rom[94][28] = 16'hFFEF;
        rom[94][29] = 16'h000C;
        rom[94][30] = 16'hFFEB;
        rom[94][31] = 16'hFFC4;
        rom[94][32] = 16'hFFF5;
        rom[94][33] = 16'hFFE1;
        rom[94][34] = 16'hFFAE;
        rom[94][35] = 16'hFFF0;
        rom[94][36] = 16'hFFF8;
        rom[94][37] = 16'hFFBB;
        rom[94][38] = 16'hFFDE;
        rom[94][39] = 16'hFFE5;
        rom[94][40] = 16'h0017;
        rom[94][41] = 16'hFFEA;
        rom[94][42] = 16'h0018;
        rom[94][43] = 16'h0010;
        rom[94][44] = 16'hFFEF;
        rom[94][45] = 16'hFFF6;
        rom[94][46] = 16'hFFDA;
        rom[94][47] = 16'hFFFB;
        rom[94][48] = 16'hFFE3;
        rom[94][49] = 16'h0033;
        rom[94][50] = 16'hFFEF;
        rom[94][51] = 16'hFFFE;
        rom[94][52] = 16'h0006;
        rom[94][53] = 16'h0010;
        rom[94][54] = 16'hFFCD;
        rom[94][55] = 16'h0033;
        rom[94][56] = 16'hFFDF;
        rom[94][57] = 16'hFFEC;
        rom[94][58] = 16'hFFF2;
        rom[94][59] = 16'hFFD7;
        rom[94][60] = 16'hFFCF;
        rom[94][61] = 16'hFFEA;
        rom[94][62] = 16'h000D;
        rom[94][63] = 16'hFFE3;
        rom[94][64] = 16'h0030;
        rom[94][65] = 16'hFFBB;
        rom[94][66] = 16'hFFCE;
        rom[94][67] = 16'h0004;
        rom[94][68] = 16'hFFF9;
        rom[94][69] = 16'h0015;
        rom[94][70] = 16'hFFFA;
        rom[94][71] = 16'h0022;
        rom[94][72] = 16'hFFB6;
        rom[94][73] = 16'hFFEF;
        rom[94][74] = 16'h0001;
        rom[94][75] = 16'hFFCC;
        rom[94][76] = 16'h0028;
        rom[94][77] = 16'hFFF1;
        rom[94][78] = 16'hFFF9;
        rom[94][79] = 16'hFFEF;
        rom[94][80] = 16'h0014;
        rom[94][81] = 16'hFFC8;
        rom[94][82] = 16'h0005;
        rom[94][83] = 16'h002D;
        rom[94][84] = 16'hFFAB;
        rom[94][85] = 16'hFFED;
        rom[94][86] = 16'hFFDF;
        rom[94][87] = 16'h0003;
        rom[94][88] = 16'hFFE6;
        rom[94][89] = 16'hFFE0;
        rom[94][90] = 16'h0009;
        rom[94][91] = 16'h0019;
        rom[94][92] = 16'h000C;
        rom[94][93] = 16'hFFF3;
        rom[94][94] = 16'hFFF4;
        rom[94][95] = 16'hFFEF;
        rom[94][96] = 16'h0001;
        rom[94][97] = 16'h0016;
        rom[94][98] = 16'hFFFD;
        rom[94][99] = 16'hFFE2;
        rom[94][100] = 16'h0017;
        rom[94][101] = 16'hFFE5;
        rom[94][102] = 16'h0025;
        rom[94][103] = 16'h001E;
        rom[94][104] = 16'hFFF9;
        rom[94][105] = 16'h000E;
        rom[94][106] = 16'hFFBF;
        rom[94][107] = 16'hFFFB;
        rom[94][108] = 16'h001B;
        rom[94][109] = 16'hFFED;
        rom[94][110] = 16'hFFD2;
        rom[94][111] = 16'h0005;
        rom[94][112] = 16'hFFE5;
        rom[94][113] = 16'h0005;
        rom[94][114] = 16'h0018;
        rom[94][115] = 16'h001B;
        rom[94][116] = 16'hFFEE;
        rom[94][117] = 16'hFFEF;
        rom[94][118] = 16'hFFDF;
        rom[94][119] = 16'hFFD7;
        rom[94][120] = 16'hFFF0;
        rom[94][121] = 16'hFFEC;
        rom[94][122] = 16'h0018;
        rom[94][123] = 16'hFFD4;
        rom[94][124] = 16'hFFE1;
        rom[94][125] = 16'hFFEB;
        rom[94][126] = 16'h0023;
        rom[94][127] = 16'hFFF8;
        rom[95][0] = 16'h001F;
        rom[95][1] = 16'hFFF6;
        rom[95][2] = 16'h0001;
        rom[95][3] = 16'hFFED;
        rom[95][4] = 16'h0022;
        rom[95][5] = 16'h000A;
        rom[95][6] = 16'h0004;
        rom[95][7] = 16'h0033;
        rom[95][8] = 16'hFFF8;
        rom[95][9] = 16'hFFEA;
        rom[95][10] = 16'hFFC8;
        rom[95][11] = 16'hFFEA;
        rom[95][12] = 16'hFFD7;
        rom[95][13] = 16'h002F;
        rom[95][14] = 16'h0006;
        rom[95][15] = 16'hFFE2;
        rom[95][16] = 16'hFFE9;
        rom[95][17] = 16'h0037;
        rom[95][18] = 16'h0007;
        rom[95][19] = 16'hFFF9;
        rom[95][20] = 16'h001B;
        rom[95][21] = 16'h001F;
        rom[95][22] = 16'hFFD9;
        rom[95][23] = 16'h0005;
        rom[95][24] = 16'h000A;
        rom[95][25] = 16'hFFF6;
        rom[95][26] = 16'h001C;
        rom[95][27] = 16'h001E;
        rom[95][28] = 16'h0018;
        rom[95][29] = 16'hFFEF;
        rom[95][30] = 16'h0010;
        rom[95][31] = 16'hFFE9;
        rom[95][32] = 16'h0012;
        rom[95][33] = 16'h0006;
        rom[95][34] = 16'h0005;
        rom[95][35] = 16'h000A;
        rom[95][36] = 16'hFFF6;
        rom[95][37] = 16'h0001;
        rom[95][38] = 16'hFFF9;
        rom[95][39] = 16'hFFFC;
        rom[95][40] = 16'hFFE8;
        rom[95][41] = 16'hFFD1;
        rom[95][42] = 16'h0003;
        rom[95][43] = 16'hFFDD;
        rom[95][44] = 16'hFFD7;
        rom[95][45] = 16'hFFDE;
        rom[95][46] = 16'hFFEE;
        rom[95][47] = 16'hFFC7;
        rom[95][48] = 16'h0012;
        rom[95][49] = 16'h0011;
        rom[95][50] = 16'hFFB1;
        rom[95][51] = 16'hFFF5;
        rom[95][52] = 16'hFFE3;
        rom[95][53] = 16'hFFE4;
        rom[95][54] = 16'hFFFA;
        rom[95][55] = 16'h0004;
        rom[95][56] = 16'h0015;
        rom[95][57] = 16'h0029;
        rom[95][58] = 16'hFFDC;
        rom[95][59] = 16'h0020;
        rom[95][60] = 16'hFFDF;
        rom[95][61] = 16'hFFF8;
        rom[95][62] = 16'hFFF9;
        rom[95][63] = 16'h0039;
        rom[95][64] = 16'hFFFA;
        rom[95][65] = 16'h001B;
        rom[95][66] = 16'h003A;
        rom[95][67] = 16'h000A;
        rom[95][68] = 16'hFFDA;
        rom[95][69] = 16'hFFCA;
        rom[95][70] = 16'hFFFA;
        rom[95][71] = 16'hFFF9;
        rom[95][72] = 16'h002E;
        rom[95][73] = 16'hFFFD;
        rom[95][74] = 16'hFFF3;
        rom[95][75] = 16'hFFDC;
        rom[95][76] = 16'hFFE3;
        rom[95][77] = 16'hFFFB;
        rom[95][78] = 16'hFFF7;
        rom[95][79] = 16'hFFE8;
        rom[95][80] = 16'h000A;
        rom[95][81] = 16'h0008;
        rom[95][82] = 16'h0004;
        rom[95][83] = 16'hFFD8;
        rom[95][84] = 16'hFFEF;
        rom[95][85] = 16'h0004;
        rom[95][86] = 16'h0009;
        rom[95][87] = 16'h001C;
        rom[95][88] = 16'h000F;
        rom[95][89] = 16'h0014;
        rom[95][90] = 16'h0024;
        rom[95][91] = 16'hFFFC;
        rom[95][92] = 16'h0010;
        rom[95][93] = 16'h0009;
        rom[95][94] = 16'hFFF0;
        rom[95][95] = 16'h0019;
        rom[95][96] = 16'hFFFA;
        rom[95][97] = 16'h001C;
        rom[95][98] = 16'hFFDD;
        rom[95][99] = 16'hFFFE;
        rom[95][100] = 16'h0006;
        rom[95][101] = 16'hFFFE;
        rom[95][102] = 16'h001A;
        rom[95][103] = 16'hFFE0;
        rom[95][104] = 16'h0011;
        rom[95][105] = 16'hFFF0;
        rom[95][106] = 16'hFFEF;
        rom[95][107] = 16'hFFCC;
        rom[95][108] = 16'h0013;
        rom[95][109] = 16'h0010;
        rom[95][110] = 16'h0011;
        rom[95][111] = 16'hFFF0;
        rom[95][112] = 16'hFFFF;
        rom[95][113] = 16'hFFF4;
        rom[95][114] = 16'h000E;
        rom[95][115] = 16'hFFEA;
        rom[95][116] = 16'hFFE7;
        rom[95][117] = 16'h000D;
        rom[95][118] = 16'h001B;
        rom[95][119] = 16'hFFDC;
        rom[95][120] = 16'h0005;
        rom[95][121] = 16'h0024;
        rom[95][122] = 16'hFFF5;
        rom[95][123] = 16'h0007;
        rom[95][124] = 16'h0001;
        rom[95][125] = 16'hFFFE;
        rom[95][126] = 16'hFFE2;
        rom[95][127] = 16'hFFD4;
        rom[96][0] = 16'h0033;
        rom[96][1] = 16'hFFE5;
        rom[96][2] = 16'hFFEE;
        rom[96][3] = 16'h0001;
        rom[96][4] = 16'h0016;
        rom[96][5] = 16'hFFE8;
        rom[96][6] = 16'hFFFC;
        rom[96][7] = 16'hFFD5;
        rom[96][8] = 16'hFFFD;
        rom[96][9] = 16'hFFC5;
        rom[96][10] = 16'h0007;
        rom[96][11] = 16'hFFD7;
        rom[96][12] = 16'hFFF4;
        rom[96][13] = 16'hFFF4;
        rom[96][14] = 16'hFFEC;
        rom[96][15] = 16'h0013;
        rom[96][16] = 16'h0039;
        rom[96][17] = 16'hFFDB;
        rom[96][18] = 16'hFFE1;
        rom[96][19] = 16'hFFF5;
        rom[96][20] = 16'hFFC5;
        rom[96][21] = 16'hFFDF;
        rom[96][22] = 16'h0003;
        rom[96][23] = 16'hFFCA;
        rom[96][24] = 16'hFFEF;
        rom[96][25] = 16'hFFB6;
        rom[96][26] = 16'hFFED;
        rom[96][27] = 16'hFFD5;
        rom[96][28] = 16'hFFF4;
        rom[96][29] = 16'hFFDA;
        rom[96][30] = 16'hFFEF;
        rom[96][31] = 16'h0025;
        rom[96][32] = 16'hFFDC;
        rom[96][33] = 16'hFFEA;
        rom[96][34] = 16'h0016;
        rom[96][35] = 16'h0007;
        rom[96][36] = 16'hFFFD;
        rom[96][37] = 16'hFFD1;
        rom[96][38] = 16'hFFE8;
        rom[96][39] = 16'h0028;
        rom[96][40] = 16'hFFF4;
        rom[96][41] = 16'hFFE7;
        rom[96][42] = 16'hFFF5;
        rom[96][43] = 16'hFFF9;
        rom[96][44] = 16'h001D;
        rom[96][45] = 16'hFFFB;
        rom[96][46] = 16'hFFE3;
        rom[96][47] = 16'h0005;
        rom[96][48] = 16'h0018;
        rom[96][49] = 16'h0005;
        rom[96][50] = 16'hFFFF;
        rom[96][51] = 16'h0031;
        rom[96][52] = 16'hFFF1;
        rom[96][53] = 16'h000C;
        rom[96][54] = 16'hFFD3;
        rom[96][55] = 16'hFFED;
        rom[96][56] = 16'hFFE0;
        rom[96][57] = 16'h0017;
        rom[96][58] = 16'h000A;
        rom[96][59] = 16'hFFD7;
        rom[96][60] = 16'h0035;
        rom[96][61] = 16'hFFF9;
        rom[96][62] = 16'hFFFE;
        rom[96][63] = 16'hFFE1;
        rom[96][64] = 16'h0016;
        rom[96][65] = 16'hFFDA;
        rom[96][66] = 16'hFFF5;
        rom[96][67] = 16'h000B;
        rom[96][68] = 16'hFFFE;
        rom[96][69] = 16'h0018;
        rom[96][70] = 16'hFFE7;
        rom[96][71] = 16'h0029;
        rom[96][72] = 16'h0007;
        rom[96][73] = 16'hFFED;
        rom[96][74] = 16'h0029;
        rom[96][75] = 16'hFFCF;
        rom[96][76] = 16'hFFD8;
        rom[96][77] = 16'h0009;
        rom[96][78] = 16'h0011;
        rom[96][79] = 16'h000C;
        rom[96][80] = 16'hFFE4;
        rom[96][81] = 16'hFFD7;
        rom[96][82] = 16'hFFE1;
        rom[96][83] = 16'hFFFD;
        rom[96][84] = 16'h000B;
        rom[96][85] = 16'h001F;
        rom[96][86] = 16'h0014;
        rom[96][87] = 16'h001B;
        rom[96][88] = 16'hFFF4;
        rom[96][89] = 16'h001F;
        rom[96][90] = 16'hFFDC;
        rom[96][91] = 16'h0015;
        rom[96][92] = 16'hFFD9;
        rom[96][93] = 16'h0024;
        rom[96][94] = 16'hFFEC;
        rom[96][95] = 16'h0006;
        rom[96][96] = 16'h0016;
        rom[96][97] = 16'hFFFD;
        rom[96][98] = 16'h0015;
        rom[96][99] = 16'h0001;
        rom[96][100] = 16'hFFF5;
        rom[96][101] = 16'h0010;
        rom[96][102] = 16'hFFE7;
        rom[96][103] = 16'h001B;
        rom[96][104] = 16'h001B;
        rom[96][105] = 16'h0010;
        rom[96][106] = 16'hFFBE;
        rom[96][107] = 16'h0023;
        rom[96][108] = 16'hFFB2;
        rom[96][109] = 16'h0009;
        rom[96][110] = 16'h0007;
        rom[96][111] = 16'h0034;
        rom[96][112] = 16'hFFB0;
        rom[96][113] = 16'hFFBB;
        rom[96][114] = 16'h000C;
        rom[96][115] = 16'hFFEB;
        rom[96][116] = 16'hFFD5;
        rom[96][117] = 16'hFFFE;
        rom[96][118] = 16'hFFCD;
        rom[96][119] = 16'hFFD5;
        rom[96][120] = 16'hFFF9;
        rom[96][121] = 16'h0026;
        rom[96][122] = 16'h0005;
        rom[96][123] = 16'hFFBF;
        rom[96][124] = 16'hFFF8;
        rom[96][125] = 16'h001E;
        rom[96][126] = 16'h0007;
        rom[96][127] = 16'h002C;
        rom[97][0] = 16'hFFFF;
        rom[97][1] = 16'hFFBF;
        rom[97][2] = 16'hFFEF;
        rom[97][3] = 16'hFFFA;
        rom[97][4] = 16'hFFDF;
        rom[97][5] = 16'hFFCB;
        rom[97][6] = 16'h0000;
        rom[97][7] = 16'hFFF1;
        rom[97][8] = 16'hFFE5;
        rom[97][9] = 16'h0010;
        rom[97][10] = 16'hFFFF;
        rom[97][11] = 16'h000B;
        rom[97][12] = 16'hFFE4;
        rom[97][13] = 16'h0041;
        rom[97][14] = 16'h001F;
        rom[97][15] = 16'hFFD6;
        rom[97][16] = 16'h0006;
        rom[97][17] = 16'h000C;
        rom[97][18] = 16'h001A;
        rom[97][19] = 16'hFFF2;
        rom[97][20] = 16'hFFFC;
        rom[97][21] = 16'hFFCD;
        rom[97][22] = 16'hFFF3;
        rom[97][23] = 16'hFFF4;
        rom[97][24] = 16'h0003;
        rom[97][25] = 16'hFFF5;
        rom[97][26] = 16'hFFFB;
        rom[97][27] = 16'h003A;
        rom[97][28] = 16'h0024;
        rom[97][29] = 16'h0012;
        rom[97][30] = 16'hFFDE;
        rom[97][31] = 16'h0027;
        rom[97][32] = 16'h001F;
        rom[97][33] = 16'h0004;
        rom[97][34] = 16'h0030;
        rom[97][35] = 16'h000D;
        rom[97][36] = 16'hFFD6;
        rom[97][37] = 16'hFFE7;
        rom[97][38] = 16'hFFFB;
        rom[97][39] = 16'h0015;
        rom[97][40] = 16'hFFC1;
        rom[97][41] = 16'hFFB4;
        rom[97][42] = 16'hFFEA;
        rom[97][43] = 16'hFFE5;
        rom[97][44] = 16'h000C;
        rom[97][45] = 16'h0000;
        rom[97][46] = 16'hFFEB;
        rom[97][47] = 16'hFFE3;
        rom[97][48] = 16'hFFC5;
        rom[97][49] = 16'hFFFB;
        rom[97][50] = 16'h0009;
        rom[97][51] = 16'h0002;
        rom[97][52] = 16'h0014;
        rom[97][53] = 16'h0000;
        rom[97][54] = 16'hFFB4;
        rom[97][55] = 16'h0017;
        rom[97][56] = 16'hFFC2;
        rom[97][57] = 16'hFFE4;
        rom[97][58] = 16'h0004;
        rom[97][59] = 16'h000A;
        rom[97][60] = 16'hFFD2;
        rom[97][61] = 16'h0024;
        rom[97][62] = 16'h002F;
        rom[97][63] = 16'hFFF9;
        rom[97][64] = 16'h0028;
        rom[97][65] = 16'hFFDE;
        rom[97][66] = 16'hFFC6;
        rom[97][67] = 16'hFFBC;
        rom[97][68] = 16'hFFD7;
        rom[97][69] = 16'hFFEA;
        rom[97][70] = 16'hFFDC;
        rom[97][71] = 16'h0013;
        rom[97][72] = 16'hFFF4;
        rom[97][73] = 16'hFFBA;
        rom[97][74] = 16'hFFF0;
        rom[97][75] = 16'hFFD2;
        rom[97][76] = 16'h0012;
        rom[97][77] = 16'hFFEF;
        rom[97][78] = 16'hFFDB;
        rom[97][79] = 16'h0008;
        rom[97][80] = 16'h0007;
        rom[97][81] = 16'hFFC5;
        rom[97][82] = 16'hFFEA;
        rom[97][83] = 16'hFFF5;
        rom[97][84] = 16'h0024;
        rom[97][85] = 16'h001B;
        rom[97][86] = 16'hFFF2;
        rom[97][87] = 16'h0026;
        rom[97][88] = 16'h0016;
        rom[97][89] = 16'hFFBD;
        rom[97][90] = 16'h000B;
        rom[97][91] = 16'h0023;
        rom[97][92] = 16'h0023;
        rom[97][93] = 16'hFFEF;
        rom[97][94] = 16'hFFF9;
        rom[97][95] = 16'hFFEA;
        rom[97][96] = 16'hFFEA;
        rom[97][97] = 16'hFFC3;
        rom[97][98] = 16'h0011;
        rom[97][99] = 16'hFFE5;
        rom[97][100] = 16'h0016;
        rom[97][101] = 16'hFFF1;
        rom[97][102] = 16'h000C;
        rom[97][103] = 16'hFFF6;
        rom[97][104] = 16'hFFF3;
        rom[97][105] = 16'hFFD6;
        rom[97][106] = 16'hFFEF;
        rom[97][107] = 16'hFFD6;
        rom[97][108] = 16'h002E;
        rom[97][109] = 16'hFFF4;
        rom[97][110] = 16'hFFF8;
        rom[97][111] = 16'hFFEF;
        rom[97][112] = 16'h0012;
        rom[97][113] = 16'h0031;
        rom[97][114] = 16'h0016;
        rom[97][115] = 16'hFFF9;
        rom[97][116] = 16'h0012;
        rom[97][117] = 16'hFFF4;
        rom[97][118] = 16'hFFEF;
        rom[97][119] = 16'hFFD4;
        rom[97][120] = 16'hFFF9;
        rom[97][121] = 16'h0016;
        rom[97][122] = 16'h0017;
        rom[97][123] = 16'h002E;
        rom[97][124] = 16'h0018;
        rom[97][125] = 16'hFFF5;
        rom[97][126] = 16'h0023;
        rom[97][127] = 16'hFFF8;
        rom[98][0] = 16'hFFE0;
        rom[98][1] = 16'hFFF9;
        rom[98][2] = 16'h001C;
        rom[98][3] = 16'h0005;
        rom[98][4] = 16'hFFE4;
        rom[98][5] = 16'h0012;
        rom[98][6] = 16'hFFC4;
        rom[98][7] = 16'h0006;
        rom[98][8] = 16'h0005;
        rom[98][9] = 16'h0030;
        rom[98][10] = 16'h0011;
        rom[98][11] = 16'hFFDC;
        rom[98][12] = 16'hFFCD;
        rom[98][13] = 16'hFFF6;
        rom[98][14] = 16'hFFF4;
        rom[98][15] = 16'h0001;
        rom[98][16] = 16'hFFC2;
        rom[98][17] = 16'h002B;
        rom[98][18] = 16'h000E;
        rom[98][19] = 16'h0035;
        rom[98][20] = 16'hFFC3;
        rom[98][21] = 16'h001A;
        rom[98][22] = 16'h002D;
        rom[98][23] = 16'h0023;
        rom[98][24] = 16'h0012;
        rom[98][25] = 16'hFFCD;
        rom[98][26] = 16'h0004;
        rom[98][27] = 16'hFFB1;
        rom[98][28] = 16'h0012;
        rom[98][29] = 16'h0006;
        rom[98][30] = 16'hFFE8;
        rom[98][31] = 16'hFFEF;
        rom[98][32] = 16'h0011;
        rom[98][33] = 16'hFFF6;
        rom[98][34] = 16'hFFBA;
        rom[98][35] = 16'h000B;
        rom[98][36] = 16'hFFE8;
        rom[98][37] = 16'hFFE7;
        rom[98][38] = 16'h001B;
        rom[98][39] = 16'hFFEC;
        rom[98][40] = 16'h000F;
        rom[98][41] = 16'h0011;
        rom[98][42] = 16'hFFDE;
        rom[98][43] = 16'h0013;
        rom[98][44] = 16'hFFE4;
        rom[98][45] = 16'h0029;
        rom[98][46] = 16'hFFFB;
        rom[98][47] = 16'hFFEF;
        rom[98][48] = 16'hFFE3;
        rom[98][49] = 16'hFFEE;
        rom[98][50] = 16'h000D;
        rom[98][51] = 16'hFFFB;
        rom[98][52] = 16'h0006;
        rom[98][53] = 16'h0007;
        rom[98][54] = 16'h000B;
        rom[98][55] = 16'hFFDF;
        rom[98][56] = 16'h0000;
        rom[98][57] = 16'hFFE9;
        rom[98][58] = 16'hFFE6;
        rom[98][59] = 16'hFFF3;
        rom[98][60] = 16'h0068;
        rom[98][61] = 16'hFFE6;
        rom[98][62] = 16'hFFE2;
        rom[98][63] = 16'h0015;
        rom[98][64] = 16'hFFFD;
        rom[98][65] = 16'hFFFA;
        rom[98][66] = 16'h0010;
        rom[98][67] = 16'hFFE9;
        rom[98][68] = 16'h0008;
        rom[98][69] = 16'hFFDF;
        rom[98][70] = 16'h002A;
        rom[98][71] = 16'h000D;
        rom[98][72] = 16'hFFE2;
        rom[98][73] = 16'h000D;
        rom[98][74] = 16'h0008;
        rom[98][75] = 16'hFFF5;
        rom[98][76] = 16'hFFEA;
        rom[98][77] = 16'hFFF7;
        rom[98][78] = 16'h0000;
        rom[98][79] = 16'hFFF6;
        rom[98][80] = 16'h0018;
        rom[98][81] = 16'hFFF0;
        rom[98][82] = 16'h0021;
        rom[98][83] = 16'hFFFD;
        rom[98][84] = 16'hFFC7;
        rom[98][85] = 16'h0001;
        rom[98][86] = 16'h0011;
        rom[98][87] = 16'hFFCD;
        rom[98][88] = 16'hFFD1;
        rom[98][89] = 16'h0006;
        rom[98][90] = 16'h000C;
        rom[98][91] = 16'hFFD7;
        rom[98][92] = 16'hFFD7;
        rom[98][93] = 16'h000C;
        rom[98][94] = 16'hFFF5;
        rom[98][95] = 16'hFFE1;
        rom[98][96] = 16'h000B;
        rom[98][97] = 16'hFFD3;
        rom[98][98] = 16'hFFE2;
        rom[98][99] = 16'hFFDA;
        rom[98][100] = 16'h002A;
        rom[98][101] = 16'hFFDF;
        rom[98][102] = 16'hFFEA;
        rom[98][103] = 16'hFFDC;
        rom[98][104] = 16'h0003;
        rom[98][105] = 16'hFFE0;
        rom[98][106] = 16'h000A;
        rom[98][107] = 16'hFFF2;
        rom[98][108] = 16'hFFD2;
        rom[98][109] = 16'h0002;
        rom[98][110] = 16'hFFFD;
        rom[98][111] = 16'hFFD6;
        rom[98][112] = 16'hFFD3;
        rom[98][113] = 16'hFFD1;
        rom[98][114] = 16'hFFC3;
        rom[98][115] = 16'hFFBC;
        rom[98][116] = 16'h000C;
        rom[98][117] = 16'h000C;
        rom[98][118] = 16'h0011;
        rom[98][119] = 16'h0000;
        rom[98][120] = 16'hFFD1;
        rom[98][121] = 16'h001F;
        rom[98][122] = 16'hFFF0;
        rom[98][123] = 16'hFFA9;
        rom[98][124] = 16'hFFE9;
        rom[98][125] = 16'hFFE5;
        rom[98][126] = 16'hFFF5;
        rom[98][127] = 16'h0016;
        rom[99][0] = 16'hFFDF;
        rom[99][1] = 16'hFFF8;
        rom[99][2] = 16'hFFFA;
        rom[99][3] = 16'hFFD2;
        rom[99][4] = 16'hFFFA;
        rom[99][5] = 16'h0023;
        rom[99][6] = 16'hFFE6;
        rom[99][7] = 16'hFFD2;
        rom[99][8] = 16'hFFFB;
        rom[99][9] = 16'hFFD7;
        rom[99][10] = 16'hFFE1;
        rom[99][11] = 16'hFFFE;
        rom[99][12] = 16'hFFDE;
        rom[99][13] = 16'hFFEF;
        rom[99][14] = 16'h0004;
        rom[99][15] = 16'h002F;
        rom[99][16] = 16'h000A;
        rom[99][17] = 16'h0018;
        rom[99][18] = 16'hFFE4;
        rom[99][19] = 16'hFFF1;
        rom[99][20] = 16'hFFB8;
        rom[99][21] = 16'hFFEF;
        rom[99][22] = 16'h001B;
        rom[99][23] = 16'hFFC3;
        rom[99][24] = 16'hFFF9;
        rom[99][25] = 16'hFFE7;
        rom[99][26] = 16'h001F;
        rom[99][27] = 16'hFFF9;
        rom[99][28] = 16'h0001;
        rom[99][29] = 16'hFFE9;
        rom[99][30] = 16'hFFFB;
        rom[99][31] = 16'hFFE5;
        rom[99][32] = 16'hFFCF;
        rom[99][33] = 16'hFFE5;
        rom[99][34] = 16'h0006;
        rom[99][35] = 16'hFFD4;
        rom[99][36] = 16'hFFCF;
        rom[99][37] = 16'h0009;
        rom[99][38] = 16'hFFE1;
        rom[99][39] = 16'hFFE4;
        rom[99][40] = 16'h0024;
        rom[99][41] = 16'hFFD5;
        rom[99][42] = 16'hFFF3;
        rom[99][43] = 16'hFFEC;
        rom[99][44] = 16'hFFDF;
        rom[99][45] = 16'h0010;
        rom[99][46] = 16'hFFB2;
        rom[99][47] = 16'hFFDC;
        rom[99][48] = 16'hFFE3;
        rom[99][49] = 16'h0016;
        rom[99][50] = 16'hFFF6;
        rom[99][51] = 16'hFFE9;
        rom[99][52] = 16'h0010;
        rom[99][53] = 16'h000B;
        rom[99][54] = 16'h001F;
        rom[99][55] = 16'hFFD7;
        rom[99][56] = 16'h0017;
        rom[99][57] = 16'hFFEA;
        rom[99][58] = 16'hFFFE;
        rom[99][59] = 16'hFFE2;
        rom[99][60] = 16'h0002;
        rom[99][61] = 16'hFFE8;
        rom[99][62] = 16'hFFDF;
        rom[99][63] = 16'hFFD3;
        rom[99][64] = 16'h0002;
        rom[99][65] = 16'hFFEB;
        rom[99][66] = 16'h0025;
        rom[99][67] = 16'h0000;
        rom[99][68] = 16'hFFEB;
        rom[99][69] = 16'h0002;
        rom[99][70] = 16'hFFF4;
        rom[99][71] = 16'h000E;
        rom[99][72] = 16'hFFEF;
        rom[99][73] = 16'h0020;
        rom[99][74] = 16'hFFCD;
        rom[99][75] = 16'hFFD9;
        rom[99][76] = 16'h0014;
        rom[99][77] = 16'h000F;
        rom[99][78] = 16'hFFE7;
        rom[99][79] = 16'hFFE2;
        rom[99][80] = 16'hFFE4;
        rom[99][81] = 16'h0006;
        rom[99][82] = 16'h000C;
        rom[99][83] = 16'hFFEA;
        rom[99][84] = 16'hFFEA;
        rom[99][85] = 16'h000B;
        rom[99][86] = 16'hFFCD;
        rom[99][87] = 16'h0024;
        rom[99][88] = 16'hFFE5;
        rom[99][89] = 16'h0016;
        rom[99][90] = 16'h0016;
        rom[99][91] = 16'h0009;
        rom[99][92] = 16'h002A;
        rom[99][93] = 16'hFFCC;
        rom[99][94] = 16'hFFF8;
        rom[99][95] = 16'hFFEA;
        rom[99][96] = 16'hFFB0;
        rom[99][97] = 16'hFFCB;
        rom[99][98] = 16'hFFFC;
        rom[99][99] = 16'h0005;
        rom[99][100] = 16'h0014;
        rom[99][101] = 16'h001F;
        rom[99][102] = 16'h001D;
        rom[99][103] = 16'hFFE2;
        rom[99][104] = 16'hFFF4;
        rom[99][105] = 16'hFFF9;
        rom[99][106] = 16'h001F;
        rom[99][107] = 16'h0018;
        rom[99][108] = 16'h0022;
        rom[99][109] = 16'h0005;
        rom[99][110] = 16'hFFF3;
        rom[99][111] = 16'hFFE7;
        rom[99][112] = 16'hFFD9;
        rom[99][113] = 16'hFFF0;
        rom[99][114] = 16'h000A;
        rom[99][115] = 16'hFFD6;
        rom[99][116] = 16'hFFE5;
        rom[99][117] = 16'hFFFA;
        rom[99][118] = 16'hFFCB;
        rom[99][119] = 16'h0009;
        rom[99][120] = 16'h0013;
        rom[99][121] = 16'hFFDB;
        rom[99][122] = 16'h0001;
        rom[99][123] = 16'h0007;
        rom[99][124] = 16'h0017;
        rom[99][125] = 16'hFFEF;
        rom[99][126] = 16'hFFF4;
        rom[99][127] = 16'hFFF0;
        rom[100][0] = 16'h000C;
        rom[100][1] = 16'hFFF6;
        rom[100][2] = 16'hFFF4;
        rom[100][3] = 16'hFFE3;
        rom[100][4] = 16'hFFF1;
        rom[100][5] = 16'hFFD3;
        rom[100][6] = 16'h0012;
        rom[100][7] = 16'hFFD8;
        rom[100][8] = 16'h0008;
        rom[100][9] = 16'hFFEB;
        rom[100][10] = 16'h0004;
        rom[100][11] = 16'hFFF8;
        rom[100][12] = 16'hFFBF;
        rom[100][13] = 16'hFFE2;
        rom[100][14] = 16'hFFEF;
        rom[100][15] = 16'hFFF4;
        rom[100][16] = 16'hFFFA;
        rom[100][17] = 16'hFFDE;
        rom[100][18] = 16'h0002;
        rom[100][19] = 16'h0012;
        rom[100][20] = 16'h0008;
        rom[100][21] = 16'h0002;
        rom[100][22] = 16'hFF9A;
        rom[100][23] = 16'hFFF2;
        rom[100][24] = 16'h001D;
        rom[100][25] = 16'h0009;
        rom[100][26] = 16'hFFEA;
        rom[100][27] = 16'h000C;
        rom[100][28] = 16'h0015;
        rom[100][29] = 16'h0009;
        rom[100][30] = 16'hFFF9;
        rom[100][31] = 16'h002E;
        rom[100][32] = 16'h001B;
        rom[100][33] = 16'hFFDF;
        rom[100][34] = 16'h001C;
        rom[100][35] = 16'h000C;
        rom[100][36] = 16'hFFF9;
        rom[100][37] = 16'h001A;
        rom[100][38] = 16'hFFD8;
        rom[100][39] = 16'h0006;
        rom[100][40] = 16'hFFF6;
        rom[100][41] = 16'h000C;
        rom[100][42] = 16'hFFD9;
        rom[100][43] = 16'hFFC1;
        rom[100][44] = 16'h0016;
        rom[100][45] = 16'hFFB8;
        rom[100][46] = 16'hFFF0;
        rom[100][47] = 16'hFFF0;
        rom[100][48] = 16'hFFD6;
        rom[100][49] = 16'h0000;
        rom[100][50] = 16'hFFED;
        rom[100][51] = 16'h0002;
        rom[100][52] = 16'hFFE1;
        rom[100][53] = 16'hFFC2;
        rom[100][54] = 16'h0002;
        rom[100][55] = 16'h0003;
        rom[100][56] = 16'hFFDA;
        rom[100][57] = 16'hFFFC;
        rom[100][58] = 16'hFFD0;
        rom[100][59] = 16'h0013;
        rom[100][60] = 16'hFFFA;
        rom[100][61] = 16'h0016;
        rom[100][62] = 16'h002F;
        rom[100][63] = 16'h0011;
        rom[100][64] = 16'h0012;
        rom[100][65] = 16'hFFD1;
        rom[100][66] = 16'hFFCB;
        rom[100][67] = 16'hFFC9;
        rom[100][68] = 16'hFFBF;
        rom[100][69] = 16'hFFE1;
        rom[100][70] = 16'hFFDB;
        rom[100][71] = 16'hFFC5;
        rom[100][72] = 16'hFFEF;
        rom[100][73] = 16'hFFEF;
        rom[100][74] = 16'h0001;
        rom[100][75] = 16'hFFDB;
        rom[100][76] = 16'hFFE2;
        rom[100][77] = 16'hFFB6;
        rom[100][78] = 16'h000D;
        rom[100][79] = 16'hFFC0;
        rom[100][80] = 16'hFFFC;
        rom[100][81] = 16'hFFE1;
        rom[100][82] = 16'hFFDB;
        rom[100][83] = 16'h0016;
        rom[100][84] = 16'hFFC0;
        rom[100][85] = 16'hFFC8;
        rom[100][86] = 16'hFFFE;
        rom[100][87] = 16'hFFCF;
        rom[100][88] = 16'h0016;
        rom[100][89] = 16'hFFD9;
        rom[100][90] = 16'h0003;
        rom[100][91] = 16'h0008;
        rom[100][92] = 16'h0005;
        rom[100][93] = 16'hFFFC;
        rom[100][94] = 16'hFFBF;
        rom[100][95] = 16'h0004;
        rom[100][96] = 16'hFFF4;
        rom[100][97] = 16'h0002;
        rom[100][98] = 16'h0016;
        rom[100][99] = 16'hFFF9;
        rom[100][100] = 16'h0020;
        rom[100][101] = 16'hFFFF;
        rom[100][102] = 16'h0006;
        rom[100][103] = 16'hFFE1;
        rom[100][104] = 16'hFFE4;
        rom[100][105] = 16'h0000;
        rom[100][106] = 16'hFFF3;
        rom[100][107] = 16'hFFE7;
        rom[100][108] = 16'h0011;
        rom[100][109] = 16'h0006;
        rom[100][110] = 16'hFFF9;
        rom[100][111] = 16'h0011;
        rom[100][112] = 16'hFFF2;
        rom[100][113] = 16'hFFFE;
        rom[100][114] = 16'h0011;
        rom[100][115] = 16'hFFFB;
        rom[100][116] = 16'hFFE1;
        rom[100][117] = 16'hFFF7;
        rom[100][118] = 16'hFFDC;
        rom[100][119] = 16'hFFD9;
        rom[100][120] = 16'hFFF0;
        rom[100][121] = 16'h0010;
        rom[100][122] = 16'hFFDC;
        rom[100][123] = 16'h0004;
        rom[100][124] = 16'hFFD4;
        rom[100][125] = 16'hFFD0;
        rom[100][126] = 16'hFFCD;
        rom[100][127] = 16'h0006;
        rom[101][0] = 16'hFFF0;
        rom[101][1] = 16'hFFC9;
        rom[101][2] = 16'hFFE8;
        rom[101][3] = 16'h000F;
        rom[101][4] = 16'h0005;
        rom[101][5] = 16'hFFEE;
        rom[101][6] = 16'hFFCF;
        rom[101][7] = 16'hFFB0;
        rom[101][8] = 16'hFFDF;
        rom[101][9] = 16'hFFD5;
        rom[101][10] = 16'h0016;
        rom[101][11] = 16'hFFF4;
        rom[101][12] = 16'h000A;
        rom[101][13] = 16'hFFFE;
        rom[101][14] = 16'hFFE1;
        rom[101][15] = 16'hFFEF;
        rom[101][16] = 16'h000E;
        rom[101][17] = 16'hFFEB;
        rom[101][18] = 16'hFFF4;
        rom[101][19] = 16'hFFF2;
        rom[101][20] = 16'hFFB7;
        rom[101][21] = 16'hFFE4;
        rom[101][22] = 16'h003A;
        rom[101][23] = 16'hFFCD;
        rom[101][24] = 16'hFFD6;
        rom[101][25] = 16'hFFCB;
        rom[101][26] = 16'h0002;
        rom[101][27] = 16'hFFF3;
        rom[101][28] = 16'h0018;
        rom[101][29] = 16'hFFCE;
        rom[101][30] = 16'h001B;
        rom[101][31] = 16'h0014;
        rom[101][32] = 16'hFFD3;
        rom[101][33] = 16'hFFEF;
        rom[101][34] = 16'hFFF6;
        rom[101][35] = 16'hFFF1;
        rom[101][36] = 16'hFFD2;
        rom[101][37] = 16'hFFF1;
        rom[101][38] = 16'hFFCD;
        rom[101][39] = 16'h0010;
        rom[101][40] = 16'h0002;
        rom[101][41] = 16'hFFBD;
        rom[101][42] = 16'h0017;
        rom[101][43] = 16'h0017;
        rom[101][44] = 16'h0027;
        rom[101][45] = 16'h0027;
        rom[101][46] = 16'hFFDA;
        rom[101][47] = 16'h002A;
        rom[101][48] = 16'hFFD2;
        rom[101][49] = 16'hFFD6;
        rom[101][50] = 16'hFFE1;
        rom[101][51] = 16'hFFFB;
        rom[101][52] = 16'h0016;
        rom[101][53] = 16'h0011;
        rom[101][54] = 16'hFFFE;
        rom[101][55] = 16'hFFE9;
        rom[101][56] = 16'h001F;
        rom[101][57] = 16'h0006;
        rom[101][58] = 16'h000E;
        rom[101][59] = 16'h0023;
        rom[101][60] = 16'h000C;
        rom[101][61] = 16'h0004;
        rom[101][62] = 16'hFFD9;
        rom[101][63] = 16'hFFD6;
        rom[101][64] = 16'h001D;
        rom[101][65] = 16'hFFD5;
        rom[101][66] = 16'hFFE7;
        rom[101][67] = 16'hFFEB;
        rom[101][68] = 16'hFFC3;
        rom[101][69] = 16'h0000;
        rom[101][70] = 16'hFFDF;
        rom[101][71] = 16'h0024;
        rom[101][72] = 16'h0013;
        rom[101][73] = 16'hFFF7;
        rom[101][74] = 16'h0024;
        rom[101][75] = 16'hFFF9;
        rom[101][76] = 16'hFFEA;
        rom[101][77] = 16'h002D;
        rom[101][78] = 16'hFFF9;
        rom[101][79] = 16'h001B;
        rom[101][80] = 16'hFFEF;
        rom[101][81] = 16'hFFF4;
        rom[101][82] = 16'hFFE7;
        rom[101][83] = 16'h002A;
        rom[101][84] = 16'hFFC0;
        rom[101][85] = 16'h0011;
        rom[101][86] = 16'hFFF6;
        rom[101][87] = 16'h000F;
        rom[101][88] = 16'hFFE0;
        rom[101][89] = 16'h001B;
        rom[101][90] = 16'hFFE7;
        rom[101][91] = 16'h0015;
        rom[101][92] = 16'hFFF4;
        rom[101][93] = 16'h001E;
        rom[101][94] = 16'hFFF0;
        rom[101][95] = 16'h002E;
        rom[101][96] = 16'h000A;
        rom[101][97] = 16'hFFD6;
        rom[101][98] = 16'h0020;
        rom[101][99] = 16'hFFE6;
        rom[101][100] = 16'h001A;
        rom[101][101] = 16'hFFFE;
        rom[101][102] = 16'hFFE1;
        rom[101][103] = 16'h0011;
        rom[101][104] = 16'h0016;
        rom[101][105] = 16'hFFCD;
        rom[101][106] = 16'hFFD4;
        rom[101][107] = 16'h0010;
        rom[101][108] = 16'hFFC3;
        rom[101][109] = 16'h0011;
        rom[101][110] = 16'h0002;
        rom[101][111] = 16'hFFF7;
        rom[101][112] = 16'h0002;
        rom[101][113] = 16'hFFED;
        rom[101][114] = 16'hFFF4;
        rom[101][115] = 16'h0006;
        rom[101][116] = 16'hFFF0;
        rom[101][117] = 16'hFFE9;
        rom[101][118] = 16'hFFF2;
        rom[101][119] = 16'hFFFA;
        rom[101][120] = 16'h0029;
        rom[101][121] = 16'h0002;
        rom[101][122] = 16'h001A;
        rom[101][123] = 16'hFFDF;
        rom[101][124] = 16'hFFFA;
        rom[101][125] = 16'h0031;
        rom[101][126] = 16'h0038;
        rom[101][127] = 16'h001F;
        rom[102][0] = 16'h000D;
        rom[102][1] = 16'h0002;
        rom[102][2] = 16'hFFE1;
        rom[102][3] = 16'hFFED;
        rom[102][4] = 16'h001F;
        rom[102][5] = 16'hFFD0;
        rom[102][6] = 16'hFFE3;
        rom[102][7] = 16'hFFFE;
        rom[102][8] = 16'hFFF7;
        rom[102][9] = 16'h001F;
        rom[102][10] = 16'hFFF1;
        rom[102][11] = 16'h0016;
        rom[102][12] = 16'h0006;
        rom[102][13] = 16'hFFE3;
        rom[102][14] = 16'hFFD5;
        rom[102][15] = 16'hFFF9;
        rom[102][16] = 16'hFFAF;
        rom[102][17] = 16'h0011;
        rom[102][18] = 16'h0007;
        rom[102][19] = 16'h0016;
        rom[102][20] = 16'h001E;
        rom[102][21] = 16'h001B;
        rom[102][22] = 16'hFFE0;
        rom[102][23] = 16'h001B;
        rom[102][24] = 16'h0013;
        rom[102][25] = 16'h0022;
        rom[102][26] = 16'h0025;
        rom[102][27] = 16'hFFE7;
        rom[102][28] = 16'h0009;
        rom[102][29] = 16'hFFE1;
        rom[102][30] = 16'h000C;
        rom[102][31] = 16'h000C;
        rom[102][32] = 16'h0006;
        rom[102][33] = 16'hFFF6;
        rom[102][34] = 16'h000F;
        rom[102][35] = 16'h000D;
        rom[102][36] = 16'hFFE9;
        rom[102][37] = 16'h0035;
        rom[102][38] = 16'h000A;
        rom[102][39] = 16'hFFDE;
        rom[102][40] = 16'hFFC8;
        rom[102][41] = 16'h0027;
        rom[102][42] = 16'hFFFE;
        rom[102][43] = 16'hFFE9;
        rom[102][44] = 16'hFFF1;
        rom[102][45] = 16'h0001;
        rom[102][46] = 16'h0014;
        rom[102][47] = 16'h0064;
        rom[102][48] = 16'hFFFE;
        rom[102][49] = 16'hFFF6;
        rom[102][50] = 16'hFFE5;
        rom[102][51] = 16'hFFD8;
        rom[102][52] = 16'hFFFD;
        rom[102][53] = 16'hFFCF;
        rom[102][54] = 16'hFFD2;
        rom[102][55] = 16'h0003;
        rom[102][56] = 16'hFFF3;
        rom[102][57] = 16'h0021;
        rom[102][58] = 16'hFFC1;
        rom[102][59] = 16'h001A;
        rom[102][60] = 16'h0010;
        rom[102][61] = 16'hFFD7;
        rom[102][62] = 16'hFFB7;
        rom[102][63] = 16'hFFF9;
        rom[102][64] = 16'hFFBA;
        rom[102][65] = 16'hFFEA;
        rom[102][66] = 16'h0018;
        rom[102][67] = 16'hFFE1;
        rom[102][68] = 16'hFFAD;
        rom[102][69] = 16'hFFD0;
        rom[102][70] = 16'h0012;
        rom[102][71] = 16'hFFF2;
        rom[102][72] = 16'h0010;
        rom[102][73] = 16'h0003;
        rom[102][74] = 16'hFFF4;
        rom[102][75] = 16'h0010;
        rom[102][76] = 16'h0011;
        rom[102][77] = 16'h0011;
        rom[102][78] = 16'hFFC3;
        rom[102][79] = 16'hFFFF;
        rom[102][80] = 16'hFFDC;
        rom[102][81] = 16'hFFF9;
        rom[102][82] = 16'h000D;
        rom[102][83] = 16'hFFF9;
        rom[102][84] = 16'hFFC1;
        rom[102][85] = 16'hFFE1;
        rom[102][86] = 16'h0001;
        rom[102][87] = 16'hFFD5;
        rom[102][88] = 16'hFFDB;
        rom[102][89] = 16'hFFF9;
        rom[102][90] = 16'h000C;
        rom[102][91] = 16'hFFB0;
        rom[102][92] = 16'h0017;
        rom[102][93] = 16'hFFD1;
        rom[102][94] = 16'hFFB5;
        rom[102][95] = 16'h000C;
        rom[102][96] = 16'hFFC4;
        rom[102][97] = 16'hFFFD;
        rom[102][98] = 16'hFFBA;
        rom[102][99] = 16'hFFFB;
        rom[102][100] = 16'hFFE7;
        rom[102][101] = 16'h0009;
        rom[102][102] = 16'hFFF7;
        rom[102][103] = 16'h0024;
        rom[102][104] = 16'hFFC8;
        rom[102][105] = 16'hFFCB;
        rom[102][106] = 16'h0002;
        rom[102][107] = 16'h0016;
        rom[102][108] = 16'hFFF9;
        rom[102][109] = 16'hFFE5;
        rom[102][110] = 16'hFFED;
        rom[102][111] = 16'hFFF7;
        rom[102][112] = 16'h000C;
        rom[102][113] = 16'hFFEB;
        rom[102][114] = 16'h0002;
        rom[102][115] = 16'h0001;
        rom[102][116] = 16'hFFF8;
        rom[102][117] = 16'h0016;
        rom[102][118] = 16'h0041;
        rom[102][119] = 16'hFFD6;
        rom[102][120] = 16'h000C;
        rom[102][121] = 16'hFFE7;
        rom[102][122] = 16'h001D;
        rom[102][123] = 16'hFFEE;
        rom[102][124] = 16'hFFDC;
        rom[102][125] = 16'hFFEE;
        rom[102][126] = 16'hFFEB;
        rom[102][127] = 16'h001F;
        rom[103][0] = 16'hFFF7;
        rom[103][1] = 16'h0019;
        rom[103][2] = 16'h0017;
        rom[103][3] = 16'hFFE9;
        rom[103][4] = 16'hFFE5;
        rom[103][5] = 16'h0013;
        rom[103][6] = 16'hFFF9;
        rom[103][7] = 16'h0035;
        rom[103][8] = 16'hFFF1;
        rom[103][9] = 16'hFFDF;
        rom[103][10] = 16'h0027;
        rom[103][11] = 16'h0002;
        rom[103][12] = 16'h0016;
        rom[103][13] = 16'hFFCC;
        rom[103][14] = 16'hFFF4;
        rom[103][15] = 16'h0019;
        rom[103][16] = 16'h000F;
        rom[103][17] = 16'hFFF1;
        rom[103][18] = 16'h0012;
        rom[103][19] = 16'h0011;
        rom[103][20] = 16'hFFF4;
        rom[103][21] = 16'hFFD9;
        rom[103][22] = 16'h0035;
        rom[103][23] = 16'hFFF5;
        rom[103][24] = 16'hFFE0;
        rom[103][25] = 16'h000E;
        rom[103][26] = 16'hFFEA;
        rom[103][27] = 16'hFFF5;
        rom[103][28] = 16'hFFD3;
        rom[103][29] = 16'h0013;
        rom[103][30] = 16'hFFE7;
        rom[103][31] = 16'hFFE4;
        rom[103][32] = 16'h0001;
        rom[103][33] = 16'h001A;
        rom[103][34] = 16'hFFF8;
        rom[103][35] = 16'h0005;
        rom[103][36] = 16'h0016;
        rom[103][37] = 16'hFFC8;
        rom[103][38] = 16'h0018;
        rom[103][39] = 16'hFFEE;
        rom[103][40] = 16'hFFFE;
        rom[103][41] = 16'hFFF9;
        rom[103][42] = 16'h0024;
        rom[103][43] = 16'hFFF0;
        rom[103][44] = 16'hFFF4;
        rom[103][45] = 16'h001F;
        rom[103][46] = 16'h002F;
        rom[103][47] = 16'h0012;
        rom[103][48] = 16'h0019;
        rom[103][49] = 16'h001B;
        rom[103][50] = 16'h0007;
        rom[103][51] = 16'hFFF9;
        rom[103][52] = 16'hFFCD;
        rom[103][53] = 16'hFFF8;
        rom[103][54] = 16'hFFE3;
        rom[103][55] = 16'hFFFA;
        rom[103][56] = 16'h0000;
        rom[103][57] = 16'h0005;
        rom[103][58] = 16'h0008;
        rom[103][59] = 16'h0019;
        rom[103][60] = 16'hFFE9;
        rom[103][61] = 16'h0046;
        rom[103][62] = 16'h0015;
        rom[103][63] = 16'h000E;
        rom[103][64] = 16'hFFF7;
        rom[103][65] = 16'hFFF9;
        rom[103][66] = 16'hFFF4;
        rom[103][67] = 16'h002A;
        rom[103][68] = 16'hFFF0;
        rom[103][69] = 16'h000E;
        rom[103][70] = 16'hFFF7;
        rom[103][71] = 16'hFFCC;
        rom[103][72] = 16'h0002;
        rom[103][73] = 16'h001B;
        rom[103][74] = 16'hFFEE;
        rom[103][75] = 16'h000C;
        rom[103][76] = 16'hFFF0;
        rom[103][77] = 16'h0014;
        rom[103][78] = 16'h000C;
        rom[103][79] = 16'h0019;
        rom[103][80] = 16'hFFF4;
        rom[103][81] = 16'h001A;
        rom[103][82] = 16'h001A;
        rom[103][83] = 16'hFFFC;
        rom[103][84] = 16'h0023;
        rom[103][85] = 16'h0002;
        rom[103][86] = 16'hFFF2;
        rom[103][87] = 16'hFFD5;
        rom[103][88] = 16'hFFE5;
        rom[103][89] = 16'h0009;
        rom[103][90] = 16'h0001;
        rom[103][91] = 16'h0005;
        rom[103][92] = 16'hFFDC;
        rom[103][93] = 16'h0022;
        rom[103][94] = 16'hFFE5;
        rom[103][95] = 16'hFFBD;
        rom[103][96] = 16'hFFEA;
        rom[103][97] = 16'hFFDB;
        rom[103][98] = 16'h0029;
        rom[103][99] = 16'h0005;
        rom[103][100] = 16'hFFCF;
        rom[103][101] = 16'hFFEC;
        rom[103][102] = 16'h001F;
        rom[103][103] = 16'hFFF2;
        rom[103][104] = 16'hFFEF;
        rom[103][105] = 16'h0017;
        rom[103][106] = 16'hFFD4;
        rom[103][107] = 16'h0007;
        rom[103][108] = 16'hFFB9;
        rom[103][109] = 16'hFFD7;
        rom[103][110] = 16'h000C;
        rom[103][111] = 16'h0001;
        rom[103][112] = 16'h0002;
        rom[103][113] = 16'hFFD9;
        rom[103][114] = 16'h0027;
        rom[103][115] = 16'hFFF9;
        rom[103][116] = 16'h001D;
        rom[103][117] = 16'hFFE9;
        rom[103][118] = 16'hFFFE;
        rom[103][119] = 16'h000A;
        rom[103][120] = 16'h0011;
        rom[103][121] = 16'hFFED;
        rom[103][122] = 16'hFFFA;
        rom[103][123] = 16'hFFEF;
        rom[103][124] = 16'hFFEB;
        rom[103][125] = 16'h000F;
        rom[103][126] = 16'hFFE5;
        rom[103][127] = 16'h001B;
        rom[104][0] = 16'hFFD3;
        rom[104][1] = 16'hFFE8;
        rom[104][2] = 16'hFFB6;
        rom[104][3] = 16'hFFEE;
        rom[104][4] = 16'h001F;
        rom[104][5] = 16'h0000;
        rom[104][6] = 16'hFFC7;
        rom[104][7] = 16'h000D;
        rom[104][8] = 16'h000C;
        rom[104][9] = 16'hFFFB;
        rom[104][10] = 16'h000E;
        rom[104][11] = 16'h001B;
        rom[104][12] = 16'hFFDA;
        rom[104][13] = 16'h0016;
        rom[104][14] = 16'hFFBC;
        rom[104][15] = 16'h0012;
        rom[104][16] = 16'hFFFA;
        rom[104][17] = 16'h0003;
        rom[104][18] = 16'h0017;
        rom[104][19] = 16'hFFDA;
        rom[104][20] = 16'h0003;
        rom[104][21] = 16'hFFEA;
        rom[104][22] = 16'h001E;
        rom[104][23] = 16'hFFEE;
        rom[104][24] = 16'h0006;
        rom[104][25] = 16'h0005;
        rom[104][26] = 16'h001A;
        rom[104][27] = 16'hFFE5;
        rom[104][28] = 16'hFFDF;
        rom[104][29] = 16'h0002;
        rom[104][30] = 16'hFFFF;
        rom[104][31] = 16'hFFF0;
        rom[104][32] = 16'h0033;
        rom[104][33] = 16'h000A;
        rom[104][34] = 16'hFFFD;
        rom[104][35] = 16'hFFF3;
        rom[104][36] = 16'hFFE7;
        rom[104][37] = 16'h0021;
        rom[104][38] = 16'hFFE7;
        rom[104][39] = 16'hFFC1;
        rom[104][40] = 16'h0011;
        rom[104][41] = 16'hFFF4;
        rom[104][42] = 16'h0011;
        rom[104][43] = 16'hFFEB;
        rom[104][44] = 16'hFFFA;
        rom[104][45] = 16'hFFFD;
        rom[104][46] = 16'h000B;
        rom[104][47] = 16'hFFDE;
        rom[104][48] = 16'h002A;
        rom[104][49] = 16'hFFDF;
        rom[104][50] = 16'hFFD8;
        rom[104][51] = 16'hFFD9;
        rom[104][52] = 16'hFFDC;
        rom[104][53] = 16'h001F;
        rom[104][54] = 16'hFFF6;
        rom[104][55] = 16'hFFDB;
        rom[104][56] = 16'h0030;
        rom[104][57] = 16'hFFCE;
        rom[104][58] = 16'hFFEF;
        rom[104][59] = 16'h002B;
        rom[104][60] = 16'h001C;
        rom[104][61] = 16'hFFF9;
        rom[104][62] = 16'hFFA3;
        rom[104][63] = 16'hFFE6;
        rom[104][64] = 16'hFFC5;
        rom[104][65] = 16'hFFD8;
        rom[104][66] = 16'hFFFE;
        rom[104][67] = 16'h0003;
        rom[104][68] = 16'hFFBF;
        rom[104][69] = 16'hFFFE;
        rom[104][70] = 16'hFFF5;
        rom[104][71] = 16'hFFE3;
        rom[104][72] = 16'h000B;
        rom[104][73] = 16'h0007;
        rom[104][74] = 16'hFFBB;
        rom[104][75] = 16'h0004;
        rom[104][76] = 16'hFFE3;
        rom[104][77] = 16'h0011;
        rom[104][78] = 16'hFFD4;
        rom[104][79] = 16'hFFF8;
        rom[104][80] = 16'hFFD2;
        rom[104][81] = 16'hFFEE;
        rom[104][82] = 16'h0018;
        rom[104][83] = 16'h0009;
        rom[104][84] = 16'h0016;
        rom[104][85] = 16'hFFF9;
        rom[104][86] = 16'hFFF4;
        rom[104][87] = 16'hFFFA;
        rom[104][88] = 16'h0011;
        rom[104][89] = 16'hFFD9;
        rom[104][90] = 16'h0037;
        rom[104][91] = 16'hFFBF;
        rom[104][92] = 16'hFFEF;
        rom[104][93] = 16'hFFCA;
        rom[104][94] = 16'h0002;
        rom[104][95] = 16'hFFD2;
        rom[104][96] = 16'hFFEA;
        rom[104][97] = 16'hFFDF;
        rom[104][98] = 16'hFFCA;
        rom[104][99] = 16'h0012;
        rom[104][100] = 16'hFFC1;
        rom[104][101] = 16'hFFF8;
        rom[104][102] = 16'hFFF2;
        rom[104][103] = 16'hFFF3;
        rom[104][104] = 16'hFFD2;
        rom[104][105] = 16'h0024;
        rom[104][106] = 16'hFFE0;
        rom[104][107] = 16'h000F;
        rom[104][108] = 16'h0002;
        rom[104][109] = 16'hFFD8;
        rom[104][110] = 16'h0003;
        rom[104][111] = 16'hFFF0;
        rom[104][112] = 16'hFFDB;
        rom[104][113] = 16'hFFB1;
        rom[104][114] = 16'hFFF2;
        rom[104][115] = 16'h000F;
        rom[104][116] = 16'hFFF6;
        rom[104][117] = 16'hFFD7;
        rom[104][118] = 16'hFFD9;
        rom[104][119] = 16'hFFC9;
        rom[104][120] = 16'h0009;
        rom[104][121] = 16'hFFBF;
        rom[104][122] = 16'h000C;
        rom[104][123] = 16'h000C;
        rom[104][124] = 16'hFFF9;
        rom[104][125] = 16'hFFFB;
        rom[104][126] = 16'hFFFC;
        rom[104][127] = 16'hFFEC;
        rom[105][0] = 16'h0017;
        rom[105][1] = 16'hFFD7;
        rom[105][2] = 16'hFFE5;
        rom[105][3] = 16'hFFC8;
        rom[105][4] = 16'hFFDD;
        rom[105][5] = 16'hFFE0;
        rom[105][6] = 16'hFFDA;
        rom[105][7] = 16'hFFF1;
        rom[105][8] = 16'hFFE1;
        rom[105][9] = 16'hFFD7;
        rom[105][10] = 16'h0024;
        rom[105][11] = 16'h0011;
        rom[105][12] = 16'hFFEF;
        rom[105][13] = 16'h0017;
        rom[105][14] = 16'h0016;
        rom[105][15] = 16'hFFE2;
        rom[105][16] = 16'h0011;
        rom[105][17] = 16'hFFFC;
        rom[105][18] = 16'hFFFC;
        rom[105][19] = 16'h000C;
        rom[105][20] = 16'h0005;
        rom[105][21] = 16'hFFDB;
        rom[105][22] = 16'hFFDB;
        rom[105][23] = 16'h0011;
        rom[105][24] = 16'hFFFE;
        rom[105][25] = 16'h0003;
        rom[105][26] = 16'h0030;
        rom[105][27] = 16'hFFFA;
        rom[105][28] = 16'h0011;
        rom[105][29] = 16'h0015;
        rom[105][30] = 16'h0029;
        rom[105][31] = 16'hFFC3;
        rom[105][32] = 16'h001B;
        rom[105][33] = 16'h0007;
        rom[105][34] = 16'hFFD2;
        rom[105][35] = 16'hFFE8;
        rom[105][36] = 16'hFFD5;
        rom[105][37] = 16'h003A;
        rom[105][38] = 16'hFFE1;
        rom[105][39] = 16'h0013;
        rom[105][40] = 16'hFFCA;
        rom[105][41] = 16'hFFFF;
        rom[105][42] = 16'hFFF1;
        rom[105][43] = 16'hFFD3;
        rom[105][44] = 16'hFFE1;
        rom[105][45] = 16'hFFEC;
        rom[105][46] = 16'hFFED;
        rom[105][47] = 16'hFF9A;
        rom[105][48] = 16'h0000;
        rom[105][49] = 16'hFFD9;
        rom[105][50] = 16'hFFC6;
        rom[105][51] = 16'h0010;
        rom[105][52] = 16'hFFE6;
        rom[105][53] = 16'h0017;
        rom[105][54] = 16'hFFAB;
        rom[105][55] = 16'hFFCF;
        rom[105][56] = 16'hFFF9;
        rom[105][57] = 16'hFFED;
        rom[105][58] = 16'hFFAA;
        rom[105][59] = 16'h0005;
        rom[105][60] = 16'hFFDC;
        rom[105][61] = 16'hFFF7;
        rom[105][62] = 16'h000A;
        rom[105][63] = 16'hFFB3;
        rom[105][64] = 16'hFFF2;
        rom[105][65] = 16'h0002;
        rom[105][66] = 16'h0002;
        rom[105][67] = 16'h0003;
        rom[105][68] = 16'hFFF2;
        rom[105][69] = 16'hFFD7;
        rom[105][70] = 16'hFFF3;
        rom[105][71] = 16'hFFE8;
        rom[105][72] = 16'hFFF7;
        rom[105][73] = 16'h000D;
        rom[105][74] = 16'hFFCE;
        rom[105][75] = 16'hFFF2;
        rom[105][76] = 16'h0002;
        rom[105][77] = 16'h0007;
        rom[105][78] = 16'h002A;
        rom[105][79] = 16'hFFDD;
        rom[105][80] = 16'hFFC8;
        rom[105][81] = 16'hFFBE;
        rom[105][82] = 16'hFFF4;
        rom[105][83] = 16'hFFFA;
        rom[105][84] = 16'hFFD7;
        rom[105][85] = 16'h0003;
        rom[105][86] = 16'h0016;
        rom[105][87] = 16'h0028;
        rom[105][88] = 16'h0005;
        rom[105][89] = 16'hFFEF;
        rom[105][90] = 16'hFFFC;
        rom[105][91] = 16'hFFF6;
        rom[105][92] = 16'hFFF9;
        rom[105][93] = 16'h0011;
        rom[105][94] = 16'hFFF7;
        rom[105][95] = 16'h0008;
        rom[105][96] = 16'h001B;
        rom[105][97] = 16'hFFF8;
        rom[105][98] = 16'hFFE2;
        rom[105][99] = 16'hFFEF;
        rom[105][100] = 16'h000D;
        rom[105][101] = 16'h001D;
        rom[105][102] = 16'hFFEA;
        rom[105][103] = 16'hFFF7;
        rom[105][104] = 16'hFFE1;
        rom[105][105] = 16'h0012;
        rom[105][106] = 16'hFFCC;
        rom[105][107] = 16'hFFE6;
        rom[105][108] = 16'h000E;
        rom[105][109] = 16'hFFF4;
        rom[105][110] = 16'hFFE4;
        rom[105][111] = 16'h0029;
        rom[105][112] = 16'h0024;
        rom[105][113] = 16'h002D;
        rom[105][114] = 16'hFFF5;
        rom[105][115] = 16'hFFEB;
        rom[105][116] = 16'h0020;
        rom[105][117] = 16'h001B;
        rom[105][118] = 16'hFFFF;
        rom[105][119] = 16'hFFBF;
        rom[105][120] = 16'h001A;
        rom[105][121] = 16'h000B;
        rom[105][122] = 16'h0016;
        rom[105][123] = 16'hFFD9;
        rom[105][124] = 16'hFFE5;
        rom[105][125] = 16'hFFE5;
        rom[105][126] = 16'hFFEE;
        rom[105][127] = 16'hFFE1;
        rom[106][0] = 16'hFFF7;
        rom[106][1] = 16'hFFD7;
        rom[106][2] = 16'h002D;
        rom[106][3] = 16'hFFFA;
        rom[106][4] = 16'h0014;
        rom[106][5] = 16'hFFA5;
        rom[106][6] = 16'hFFFF;
        rom[106][7] = 16'hFFBA;
        rom[106][8] = 16'hFFEF;
        rom[106][9] = 16'h001A;
        rom[106][10] = 16'h000E;
        rom[106][11] = 16'h0025;
        rom[106][12] = 16'hFFF4;
        rom[106][13] = 16'h001D;
        rom[106][14] = 16'hFFD9;
        rom[106][15] = 16'h001F;
        rom[106][16] = 16'h0013;
        rom[106][17] = 16'h000F;
        rom[106][18] = 16'h0017;
        rom[106][19] = 16'hFFE6;
        rom[106][20] = 16'h0016;
        rom[106][21] = 16'hFFE1;
        rom[106][22] = 16'hFFE1;
        rom[106][23] = 16'hFFEA;
        rom[106][24] = 16'h001C;
        rom[106][25] = 16'hFFF5;
        rom[106][26] = 16'hFFCD;
        rom[106][27] = 16'h000E;
        rom[106][28] = 16'hFFE2;
        rom[106][29] = 16'h0028;
        rom[106][30] = 16'hFFF7;
        rom[106][31] = 16'hFFE5;
        rom[106][32] = 16'hFFF4;
        rom[106][33] = 16'hFFF0;
        rom[106][34] = 16'hFFFF;
        rom[106][35] = 16'hFFF7;
        rom[106][36] = 16'hFFEC;
        rom[106][37] = 16'hFFF7;
        rom[106][38] = 16'h000C;
        rom[106][39] = 16'hFFDE;
        rom[106][40] = 16'h000F;
        rom[106][41] = 16'hFFF1;
        rom[106][42] = 16'hFFEA;
        rom[106][43] = 16'hFFE9;
        rom[106][44] = 16'h0002;
        rom[106][45] = 16'h0025;
        rom[106][46] = 16'h0002;
        rom[106][47] = 16'hFFBC;
        rom[106][48] = 16'hFFF1;
        rom[106][49] = 16'hFFB8;
        rom[106][50] = 16'h001C;
        rom[106][51] = 16'hFFDD;
        rom[106][52] = 16'h000E;
        rom[106][53] = 16'h0018;
        rom[106][54] = 16'h0020;
        rom[106][55] = 16'h0002;
        rom[106][56] = 16'h001B;
        rom[106][57] = 16'hFFDF;
        rom[106][58] = 16'hFFE4;
        rom[106][59] = 16'h0000;
        rom[106][60] = 16'h000C;
        rom[106][61] = 16'hFFF4;
        rom[106][62] = 16'hFFF4;
        rom[106][63] = 16'hFFB0;
        rom[106][64] = 16'h0014;
        rom[106][65] = 16'hFFF4;
        rom[106][66] = 16'h0007;
        rom[106][67] = 16'hFFD0;
        rom[106][68] = 16'hFFCF;
        rom[106][69] = 16'hFFC9;
        rom[106][70] = 16'h000C;
        rom[106][71] = 16'hFFF1;
        rom[106][72] = 16'h000C;
        rom[106][73] = 16'h0010;
        rom[106][74] = 16'hFFF4;
        rom[106][75] = 16'hFFEF;
        rom[106][76] = 16'h0003;
        rom[106][77] = 16'hFFEF;
        rom[106][78] = 16'hFFD9;
        rom[106][79] = 16'hFFF8;
        rom[106][80] = 16'hFFE0;
        rom[106][81] = 16'hFFCC;
        rom[106][82] = 16'hFF9F;
        rom[106][83] = 16'h0018;
        rom[106][84] = 16'hFFF8;
        rom[106][85] = 16'hFFF5;
        rom[106][86] = 16'h0005;
        rom[106][87] = 16'hFFFC;
        rom[106][88] = 16'hFFFE;
        rom[106][89] = 16'h0020;
        rom[106][90] = 16'hFFDC;
        rom[106][91] = 16'h001B;
        rom[106][92] = 16'h001B;
        rom[106][93] = 16'hFFDC;
        rom[106][94] = 16'h0015;
        rom[106][95] = 16'hFFEB;
        rom[106][96] = 16'hFFE8;
        rom[106][97] = 16'h0000;
        rom[106][98] = 16'hFFEF;
        rom[106][99] = 16'hFFD2;
        rom[106][100] = 16'hFFFD;
        rom[106][101] = 16'hFFFC;
        rom[106][102] = 16'h001C;
        rom[106][103] = 16'h0017;
        rom[106][104] = 16'hFFC8;
        rom[106][105] = 16'hFFE4;
        rom[106][106] = 16'h003D;
        rom[106][107] = 16'hFFFD;
        rom[106][108] = 16'h0001;
        rom[106][109] = 16'hFFD1;
        rom[106][110] = 16'hFFF2;
        rom[106][111] = 16'hFFCE;
        rom[106][112] = 16'hFFDF;
        rom[106][113] = 16'h0009;
        rom[106][114] = 16'h0013;
        rom[106][115] = 16'h0011;
        rom[106][116] = 16'hFFFD;
        rom[106][117] = 16'hFFEA;
        rom[106][118] = 16'hFFDC;
        rom[106][119] = 16'h0000;
        rom[106][120] = 16'h0029;
        rom[106][121] = 16'h0001;
        rom[106][122] = 16'h0014;
        rom[106][123] = 16'h0017;
        rom[106][124] = 16'h0020;
        rom[106][125] = 16'hFFE2;
        rom[106][126] = 16'h0008;
        rom[106][127] = 16'hFFF7;
        rom[107][0] = 16'hFFC8;
        rom[107][1] = 16'hFFE6;
        rom[107][2] = 16'h0001;
        rom[107][3] = 16'hFFCB;
        rom[107][4] = 16'h0019;
        rom[107][5] = 16'h0009;
        rom[107][6] = 16'h0018;
        rom[107][7] = 16'hFFFF;
        rom[107][8] = 16'h0024;
        rom[107][9] = 16'hFFD5;
        rom[107][10] = 16'h0029;
        rom[107][11] = 16'hFFA0;
        rom[107][12] = 16'h001B;
        rom[107][13] = 16'hFFEA;
        rom[107][14] = 16'h000E;
        rom[107][15] = 16'hFFF0;
        rom[107][16] = 16'h0038;
        rom[107][17] = 16'h0023;
        rom[107][18] = 16'hFFC8;
        rom[107][19] = 16'h0029;
        rom[107][20] = 16'hFFB8;
        rom[107][21] = 16'h0016;
        rom[107][22] = 16'hFFEF;
        rom[107][23] = 16'hFFD4;
        rom[107][24] = 16'hFFDD;
        rom[107][25] = 16'hFFB0;
        rom[107][26] = 16'h003D;
        rom[107][27] = 16'hFFBA;
        rom[107][28] = 16'hFFDB;
        rom[107][29] = 16'h0026;
        rom[107][30] = 16'h0002;
        rom[107][31] = 16'hFFF0;
        rom[107][32] = 16'hFFD8;
        rom[107][33] = 16'h002A;
        rom[107][34] = 16'hFFDD;
        rom[107][35] = 16'hFFF9;
        rom[107][36] = 16'h001B;
        rom[107][37] = 16'h0037;
        rom[107][38] = 16'hFFD5;
        rom[107][39] = 16'hFFF9;
        rom[107][40] = 16'h0016;
        rom[107][41] = 16'h0007;
        rom[107][42] = 16'h001B;
        rom[107][43] = 16'hFFE6;
        rom[107][44] = 16'h0000;
        rom[107][45] = 16'h000C;
        rom[107][46] = 16'h0020;
        rom[107][47] = 16'hFFFB;
        rom[107][48] = 16'h0001;
        rom[107][49] = 16'h0007;
        rom[107][50] = 16'hFFF4;
        rom[107][51] = 16'h001A;
        rom[107][52] = 16'h001B;
        rom[107][53] = 16'h001F;
        rom[107][54] = 16'hFFEC;
        rom[107][55] = 16'hFFD7;
        rom[107][56] = 16'h0044;
        rom[107][57] = 16'hFFF9;
        rom[107][58] = 16'h003D;
        rom[107][59] = 16'h0005;
        rom[107][60] = 16'hFFF5;
        rom[107][61] = 16'hFFFD;
        rom[107][62] = 16'hFFFC;
        rom[107][63] = 16'h0024;
        rom[107][64] = 16'hFFFE;
        rom[107][65] = 16'hFFF3;
        rom[107][66] = 16'h0018;
        rom[107][67] = 16'h0006;
        rom[107][68] = 16'h000C;
        rom[107][69] = 16'hFFAE;
        rom[107][70] = 16'hFFFA;
        rom[107][71] = 16'h001E;
        rom[107][72] = 16'hFFD8;
        rom[107][73] = 16'h0013;
        rom[107][74] = 16'h0008;
        rom[107][75] = 16'h000C;
        rom[107][76] = 16'h0029;
        rom[107][77] = 16'h0030;
        rom[107][78] = 16'hFFEE;
        rom[107][79] = 16'h0029;
        rom[107][80] = 16'h0002;
        rom[107][81] = 16'hFFEA;
        rom[107][82] = 16'h001B;
        rom[107][83] = 16'h0020;
        rom[107][84] = 16'hFFF9;
        rom[107][85] = 16'h001E;
        rom[107][86] = 16'hFFE9;
        rom[107][87] = 16'h0030;
        rom[107][88] = 16'hFFEC;
        rom[107][89] = 16'h002B;
        rom[107][90] = 16'h001B;
        rom[107][91] = 16'h0023;
        rom[107][92] = 16'h0038;
        rom[107][93] = 16'hFFDC;
        rom[107][94] = 16'hFFED;
        rom[107][95] = 16'hFFE4;
        rom[107][96] = 16'h0003;
        rom[107][97] = 16'h0037;
        rom[107][98] = 16'h0033;
        rom[107][99] = 16'h0005;
        rom[107][100] = 16'h0015;
        rom[107][101] = 16'hFFFB;
        rom[107][102] = 16'h0016;
        rom[107][103] = 16'hFFDE;
        rom[107][104] = 16'h0043;
        rom[107][105] = 16'h001B;
        rom[107][106] = 16'h001B;
        rom[107][107] = 16'hFFEF;
        rom[107][108] = 16'h0007;
        rom[107][109] = 16'hFFE1;
        rom[107][110] = 16'hFFF4;
        rom[107][111] = 16'hFFF1;
        rom[107][112] = 16'hFFAE;
        rom[107][113] = 16'h000E;
        rom[107][114] = 16'hFFF8;
        rom[107][115] = 16'hFFEA;
        rom[107][116] = 16'hFFF1;
        rom[107][117] = 16'h001C;
        rom[107][118] = 16'hFFFD;
        rom[107][119] = 16'hFFED;
        rom[107][120] = 16'hFFC3;
        rom[107][121] = 16'hFFE1;
        rom[107][122] = 16'h001B;
        rom[107][123] = 16'hFFF3;
        rom[107][124] = 16'h0000;
        rom[107][125] = 16'h001A;
        rom[107][126] = 16'hFFFF;
        rom[107][127] = 16'h0009;
        rom[108][0] = 16'hFFF9;
        rom[108][1] = 16'h0010;
        rom[108][2] = 16'h0000;
        rom[108][3] = 16'h0007;
        rom[108][4] = 16'hFFB1;
        rom[108][5] = 16'hFFF3;
        rom[108][6] = 16'hFFF4;
        rom[108][7] = 16'h0012;
        rom[108][8] = 16'hFFEF;
        rom[108][9] = 16'h0029;
        rom[108][10] = 16'h000A;
        rom[108][11] = 16'h0037;
        rom[108][12] = 16'hFFEC;
        rom[108][13] = 16'hFFFC;
        rom[108][14] = 16'hFFE0;
        rom[108][15] = 16'hFFF7;
        rom[108][16] = 16'h0000;
        rom[108][17] = 16'h0016;
        rom[108][18] = 16'h001C;
        rom[108][19] = 16'h0016;
        rom[108][20] = 16'hFFB9;
        rom[108][21] = 16'h0009;
        rom[108][22] = 16'hFFFB;
        rom[108][23] = 16'hFFE9;
        rom[108][24] = 16'hFFF9;
        rom[108][25] = 16'hFF9E;
        rom[108][26] = 16'h0015;
        rom[108][27] = 16'hFFCD;
        rom[108][28] = 16'hFFFE;
        rom[108][29] = 16'h0030;
        rom[108][30] = 16'hFFF7;
        rom[108][31] = 16'hFFE1;
        rom[108][32] = 16'h000D;
        rom[108][33] = 16'hFFEC;
        rom[108][34] = 16'hFFC9;
        rom[108][35] = 16'h0002;
        rom[108][36] = 16'h0016;
        rom[108][37] = 16'hFFD5;
        rom[108][38] = 16'h0015;
        rom[108][39] = 16'h0023;
        rom[108][40] = 16'h0024;
        rom[108][41] = 16'h0016;
        rom[108][42] = 16'h0011;
        rom[108][43] = 16'h0013;
        rom[108][44] = 16'h0003;
        rom[108][45] = 16'h0019;
        rom[108][46] = 16'h0005;
        rom[108][47] = 16'hFFCE;
        rom[108][48] = 16'h0022;
        rom[108][49] = 16'h0007;
        rom[108][50] = 16'h0000;
        rom[108][51] = 16'hFFD4;
        rom[108][52] = 16'h0015;
        rom[108][53] = 16'h0037;
        rom[108][54] = 16'h0007;
        rom[108][55] = 16'hFFDC;
        rom[108][56] = 16'hFFE5;
        rom[108][57] = 16'hFFD3;
        rom[108][58] = 16'hFFD8;
        rom[108][59] = 16'h0005;
        rom[108][60] = 16'hFFF0;
        rom[108][61] = 16'h0013;
        rom[108][62] = 16'hFFEE;
        rom[108][63] = 16'h0007;
        rom[108][64] = 16'hFFE3;
        rom[108][65] = 16'hFFF6;
        rom[108][66] = 16'hFFF4;
        rom[108][67] = 16'hFFF0;
        rom[108][68] = 16'h0011;
        rom[108][69] = 16'h0023;
        rom[108][70] = 16'h0005;
        rom[108][71] = 16'h001B;
        rom[108][72] = 16'h000E;
        rom[108][73] = 16'h0004;
        rom[108][74] = 16'hFFE3;
        rom[108][75] = 16'hFFEF;
        rom[108][76] = 16'hFFD1;
        rom[108][77] = 16'hFFE1;
        rom[108][78] = 16'h0013;
        rom[108][79] = 16'h0018;
        rom[108][80] = 16'hFFDE;
        rom[108][81] = 16'h0012;
        rom[108][82] = 16'hFFE5;
        rom[108][83] = 16'h0007;
        rom[108][84] = 16'hFFDF;
        rom[108][85] = 16'h0003;
        rom[108][86] = 16'h0002;
        rom[108][87] = 16'hFFEF;
        rom[108][88] = 16'hFFC1;
        rom[108][89] = 16'hFFFE;
        rom[108][90] = 16'hFFEA;
        rom[108][91] = 16'hFFF5;
        rom[108][92] = 16'hFFEA;
        rom[108][93] = 16'h004F;
        rom[108][94] = 16'h000C;
        rom[108][95] = 16'hFFD6;
        rom[108][96] = 16'h0027;
        rom[108][97] = 16'hFFFD;
        rom[108][98] = 16'h0002;
        rom[108][99] = 16'h0028;
        rom[108][100] = 16'h0001;
        rom[108][101] = 16'hFFC3;
        rom[108][102] = 16'hFFA2;
        rom[108][103] = 16'hFFC6;
        rom[108][104] = 16'hFFEE;
        rom[108][105] = 16'hFFDC;
        rom[108][106] = 16'hFFC3;
        rom[108][107] = 16'h002D;
        rom[108][108] = 16'hFFDE;
        rom[108][109] = 16'h0024;
        rom[108][110] = 16'hFFD3;
        rom[108][111] = 16'h0013;
        rom[108][112] = 16'h000B;
        rom[108][113] = 16'hFFDB;
        rom[108][114] = 16'h000E;
        rom[108][115] = 16'hFFF7;
        rom[108][116] = 16'hFFC0;
        rom[108][117] = 16'hFFF4;
        rom[108][118] = 16'hFFC2;
        rom[108][119] = 16'h0018;
        rom[108][120] = 16'h0025;
        rom[108][121] = 16'hFFF3;
        rom[108][122] = 16'h0011;
        rom[108][123] = 16'hFFAF;
        rom[108][124] = 16'hFFF8;
        rom[108][125] = 16'h0009;
        rom[108][126] = 16'h0009;
        rom[108][127] = 16'h003B;
        rom[109][0] = 16'h0034;
        rom[109][1] = 16'hFFCD;
        rom[109][2] = 16'h0007;
        rom[109][3] = 16'h0006;
        rom[109][4] = 16'h0001;
        rom[109][5] = 16'h0016;
        rom[109][6] = 16'hFFF8;
        rom[109][7] = 16'hFFCF;
        rom[109][8] = 16'h0021;
        rom[109][9] = 16'h0007;
        rom[109][10] = 16'hFFFE;
        rom[109][11] = 16'hFFE3;
        rom[109][12] = 16'h0011;
        rom[109][13] = 16'h000A;
        rom[109][14] = 16'hFFFA;
        rom[109][15] = 16'hFFFA;
        rom[109][16] = 16'hFFEF;
        rom[109][17] = 16'hFFE5;
        rom[109][18] = 16'hFFFF;
        rom[109][19] = 16'hFFE3;
        rom[109][20] = 16'hFFD0;
        rom[109][21] = 16'hFFFD;
        rom[109][22] = 16'h001B;
        rom[109][23] = 16'hFFE9;
        rom[109][24] = 16'h0034;
        rom[109][25] = 16'hFFDA;
        rom[109][26] = 16'hFFF3;
        rom[109][27] = 16'hFFF4;
        rom[109][28] = 16'hFFED;
        rom[109][29] = 16'hFFF5;
        rom[109][30] = 16'hFFF9;
        rom[109][31] = 16'h000B;
        rom[109][32] = 16'h001E;
        rom[109][33] = 16'h0008;
        rom[109][34] = 16'hFFC0;
        rom[109][35] = 16'h0006;
        rom[109][36] = 16'hFFEF;
        rom[109][37] = 16'hFFB1;
        rom[109][38] = 16'h002D;
        rom[109][39] = 16'h0002;
        rom[109][40] = 16'h0007;
        rom[109][41] = 16'hFFF4;
        rom[109][42] = 16'h001D;
        rom[109][43] = 16'hFFC8;
        rom[109][44] = 16'h0011;
        rom[109][45] = 16'h0011;
        rom[109][46] = 16'hFFD2;
        rom[109][47] = 16'h0002;
        rom[109][48] = 16'h0010;
        rom[109][49] = 16'h0013;
        rom[109][50] = 16'h0029;
        rom[109][51] = 16'h0038;
        rom[109][52] = 16'hFFF5;
        rom[109][53] = 16'h001B;
        rom[109][54] = 16'hFFF9;
        rom[109][55] = 16'hFFE5;
        rom[109][56] = 16'h000C;
        rom[109][57] = 16'h0006;
        rom[109][58] = 16'h000D;
        rom[109][59] = 16'hFFEE;
        rom[109][60] = 16'hFFD3;
        rom[109][61] = 16'h0003;
        rom[109][62] = 16'hFFE9;
        rom[109][63] = 16'hFFCF;
        rom[109][64] = 16'h0007;
        rom[109][65] = 16'hFFE3;
        rom[109][66] = 16'h0005;
        rom[109][67] = 16'h0011;
        rom[109][68] = 16'h0002;
        rom[109][69] = 16'hFFF9;
        rom[109][70] = 16'h0022;
        rom[109][71] = 16'h0015;
        rom[109][72] = 16'h0013;
        rom[109][73] = 16'h0000;
        rom[109][74] = 16'hFFED;
        rom[109][75] = 16'h001A;
        rom[109][76] = 16'hFFA3;
        rom[109][77] = 16'h0002;
        rom[109][78] = 16'h0036;
        rom[109][79] = 16'h0026;
        rom[109][80] = 16'hFFDF;
        rom[109][81] = 16'hFFF8;
        rom[109][82] = 16'hFFD4;
        rom[109][83] = 16'h002B;
        rom[109][84] = 16'hFFFC;
        rom[109][85] = 16'hFFD2;
        rom[109][86] = 16'hFFEC;
        rom[109][87] = 16'h000C;
        rom[109][88] = 16'hFFFD;
        rom[109][89] = 16'h0025;
        rom[109][90] = 16'hFFCD;
        rom[109][91] = 16'h0011;
        rom[109][92] = 16'hFFE1;
        rom[109][93] = 16'h0041;
        rom[109][94] = 16'hFFAC;
        rom[109][95] = 16'h0030;
        rom[109][96] = 16'h000D;
        rom[109][97] = 16'h0041;
        rom[109][98] = 16'h0009;
        rom[109][99] = 16'hFFD6;
        rom[109][100] = 16'h0014;
        rom[109][101] = 16'h000F;
        rom[109][102] = 16'hFFEA;
        rom[109][103] = 16'h0026;
        rom[109][104] = 16'h0036;
        rom[109][105] = 16'hFFD0;
        rom[109][106] = 16'hFFF4;
        rom[109][107] = 16'h0024;
        rom[109][108] = 16'hFFA1;
        rom[109][109] = 16'h001D;
        rom[109][110] = 16'h0017;
        rom[109][111] = 16'hFFE1;
        rom[109][112] = 16'hFFDB;
        rom[109][113] = 16'h0003;
        rom[109][114] = 16'h002C;
        rom[109][115] = 16'hFFE6;
        rom[109][116] = 16'hFFE2;
        rom[109][117] = 16'hFFFE;
        rom[109][118] = 16'hFFDE;
        rom[109][119] = 16'h0001;
        rom[109][120] = 16'h0033;
        rom[109][121] = 16'hFFF4;
        rom[109][122] = 16'h000C;
        rom[109][123] = 16'hFFD3;
        rom[109][124] = 16'h0027;
        rom[109][125] = 16'h0030;
        rom[109][126] = 16'h001A;
        rom[109][127] = 16'h0007;
        rom[110][0] = 16'h0032;
        rom[110][1] = 16'hFFF3;
        rom[110][2] = 16'hFFEF;
        rom[110][3] = 16'hFFFB;
        rom[110][4] = 16'h000E;
        rom[110][5] = 16'h0007;
        rom[110][6] = 16'hFFCB;
        rom[110][7] = 16'hFFD7;
        rom[110][8] = 16'h0046;
        rom[110][9] = 16'h001F;
        rom[110][10] = 16'hFFE0;
        rom[110][11] = 16'h001F;
        rom[110][12] = 16'hFFE2;
        rom[110][13] = 16'h0019;
        rom[110][14] = 16'hFFF6;
        rom[110][15] = 16'h0002;
        rom[110][16] = 16'hFFEC;
        rom[110][17] = 16'hFFEF;
        rom[110][18] = 16'hFFFE;
        rom[110][19] = 16'h0012;
        rom[110][20] = 16'hFFEF;
        rom[110][21] = 16'h0013;
        rom[110][22] = 16'hFFDA;
        rom[110][23] = 16'h0014;
        rom[110][24] = 16'h0012;
        rom[110][25] = 16'hFFF4;
        rom[110][26] = 16'hFFD9;
        rom[110][27] = 16'hFFEC;
        rom[110][28] = 16'h000A;
        rom[110][29] = 16'hFFE5;
        rom[110][30] = 16'h0004;
        rom[110][31] = 16'h0014;
        rom[110][32] = 16'hFFE2;
        rom[110][33] = 16'hFFF9;
        rom[110][34] = 16'h001B;
        rom[110][35] = 16'h000D;
        rom[110][36] = 16'hFFE4;
        rom[110][37] = 16'h000D;
        rom[110][38] = 16'h0013;
        rom[110][39] = 16'hFFF6;
        rom[110][40] = 16'h0000;
        rom[110][41] = 16'h0044;
        rom[110][42] = 16'hFFD0;
        rom[110][43] = 16'hFFF0;
        rom[110][44] = 16'hFFE3;
        rom[110][45] = 16'hFFDF;
        rom[110][46] = 16'hFFFF;
        rom[110][47] = 16'hFFEA;
        rom[110][48] = 16'hFFEE;
        rom[110][49] = 16'hFFF4;
        rom[110][50] = 16'hFFDF;
        rom[110][51] = 16'h0011;
        rom[110][52] = 16'hFFE9;
        rom[110][53] = 16'hFFE2;
        rom[110][54] = 16'hFFFF;
        rom[110][55] = 16'hFFBE;
        rom[110][56] = 16'hFFFD;
        rom[110][57] = 16'h0016;
        rom[110][58] = 16'h0006;
        rom[110][59] = 16'hFFEC;
        rom[110][60] = 16'h003F;
        rom[110][61] = 16'h001B;
        rom[110][62] = 16'hFFF9;
        rom[110][63] = 16'hFFE3;
        rom[110][64] = 16'h0006;
        rom[110][65] = 16'h001B;
        rom[110][66] = 16'h0009;
        rom[110][67] = 16'hFFFD;
        rom[110][68] = 16'h0016;
        rom[110][69] = 16'hFFD7;
        rom[110][70] = 16'h0013;
        rom[110][71] = 16'hFFC8;
        rom[110][72] = 16'h003B;
        rom[110][73] = 16'h001B;
        rom[110][74] = 16'h001D;
        rom[110][75] = 16'h0016;
        rom[110][76] = 16'h0022;
        rom[110][77] = 16'h0007;
        rom[110][78] = 16'h0003;
        rom[110][79] = 16'hFFF7;
        rom[110][80] = 16'hFFD3;
        rom[110][81] = 16'hFFD0;
        rom[110][82] = 16'hFFCD;
        rom[110][83] = 16'h001B;
        rom[110][84] = 16'hFFE8;
        rom[110][85] = 16'hFFF6;
        rom[110][86] = 16'h0025;
        rom[110][87] = 16'h001A;
        rom[110][88] = 16'h0018;
        rom[110][89] = 16'h002A;
        rom[110][90] = 16'hFFE0;
        rom[110][91] = 16'hFFD5;
        rom[110][92] = 16'h003D;
        rom[110][93] = 16'h0029;
        rom[110][94] = 16'h001F;
        rom[110][95] = 16'h0005;
        rom[110][96] = 16'h0016;
        rom[110][97] = 16'h0005;
        rom[110][98] = 16'h0000;
        rom[110][99] = 16'hFFF3;
        rom[110][100] = 16'hFFEB;
        rom[110][101] = 16'hFFFC;
        rom[110][102] = 16'hFFC3;
        rom[110][103] = 16'h000C;
        rom[110][104] = 16'h0003;
        rom[110][105] = 16'h000E;
        rom[110][106] = 16'hFFD2;
        rom[110][107] = 16'hFFFD;
        rom[110][108] = 16'hFFAC;
        rom[110][109] = 16'hFFFE;
        rom[110][110] = 16'hFFF4;
        rom[110][111] = 16'hFFFC;
        rom[110][112] = 16'hFFE5;
        rom[110][113] = 16'hFFC7;
        rom[110][114] = 16'hFFED;
        rom[110][115] = 16'hFFC4;
        rom[110][116] = 16'h0010;
        rom[110][117] = 16'h001B;
        rom[110][118] = 16'hFFEC;
        rom[110][119] = 16'hFFF5;
        rom[110][120] = 16'h0035;
        rom[110][121] = 16'hFFF5;
        rom[110][122] = 16'h0020;
        rom[110][123] = 16'h001F;
        rom[110][124] = 16'h0005;
        rom[110][125] = 16'h0008;
        rom[110][126] = 16'hFFD2;
        rom[110][127] = 16'hFFE2;
        rom[111][0] = 16'hFFF1;
        rom[111][1] = 16'h001A;
        rom[111][2] = 16'h0007;
        rom[111][3] = 16'hFFB2;
        rom[111][4] = 16'h0023;
        rom[111][5] = 16'h001F;
        rom[111][6] = 16'h0014;
        rom[111][7] = 16'h0004;
        rom[111][8] = 16'h0002;
        rom[111][9] = 16'hFFD7;
        rom[111][10] = 16'h0029;
        rom[111][11] = 16'hFFF3;
        rom[111][12] = 16'hFFFF;
        rom[111][13] = 16'hFFC3;
        rom[111][14] = 16'h0017;
        rom[111][15] = 16'h0015;
        rom[111][16] = 16'h000C;
        rom[111][17] = 16'hFFC5;
        rom[111][18] = 16'hFFE3;
        rom[111][19] = 16'h0011;
        rom[111][20] = 16'hFFF7;
        rom[111][21] = 16'hFFF4;
        rom[111][22] = 16'h000D;
        rom[111][23] = 16'hFFC8;
        rom[111][24] = 16'hFFEF;
        rom[111][25] = 16'hFFF3;
        rom[111][26] = 16'hFFF6;
        rom[111][27] = 16'h0012;
        rom[111][28] = 16'h0010;
        rom[111][29] = 16'hFFED;
        rom[111][30] = 16'hFFF8;
        rom[111][31] = 16'hFFC3;
        rom[111][32] = 16'h0007;
        rom[111][33] = 16'hFFD9;
        rom[111][34] = 16'hFFD7;
        rom[111][35] = 16'hFFE4;
        rom[111][36] = 16'h000C;
        rom[111][37] = 16'h0003;
        rom[111][38] = 16'hFFDC;
        rom[111][39] = 16'hFFFE;
        rom[111][40] = 16'hFFE0;
        rom[111][41] = 16'hFFEE;
        rom[111][42] = 16'hFFF4;
        rom[111][43] = 16'hFFD3;
        rom[111][44] = 16'hFFEA;
        rom[111][45] = 16'hFFE6;
        rom[111][46] = 16'hFFF8;
        rom[111][47] = 16'h001F;
        rom[111][48] = 16'h000C;
        rom[111][49] = 16'h001E;
        rom[111][50] = 16'h0001;
        rom[111][51] = 16'hFFEA;
        rom[111][52] = 16'h002F;
        rom[111][53] = 16'hFFE5;
        rom[111][54] = 16'h0019;
        rom[111][55] = 16'hFFD6;
        rom[111][56] = 16'h001D;
        rom[111][57] = 16'hFFE3;
        rom[111][58] = 16'hFFDF;
        rom[111][59] = 16'hFFE0;
        rom[111][60] = 16'hFFF7;
        rom[111][61] = 16'hFFF2;
        rom[111][62] = 16'h001B;
        rom[111][63] = 16'hFFDE;
        rom[111][64] = 16'h0001;
        rom[111][65] = 16'hFFEA;
        rom[111][66] = 16'h0032;
        rom[111][67] = 16'h000E;
        rom[111][68] = 16'hFFDD;
        rom[111][69] = 16'hFFFE;
        rom[111][70] = 16'h001F;
        rom[111][71] = 16'hFFF8;
        rom[111][72] = 16'hFFDF;
        rom[111][73] = 16'h0044;
        rom[111][74] = 16'hFFE5;
        rom[111][75] = 16'hFFD2;
        rom[111][76] = 16'h0023;
        rom[111][77] = 16'h0011;
        rom[111][78] = 16'h0006;
        rom[111][79] = 16'hFFEA;
        rom[111][80] = 16'hFFF1;
        rom[111][81] = 16'h0035;
        rom[111][82] = 16'hFFEF;
        rom[111][83] = 16'h0007;
        rom[111][84] = 16'h0019;
        rom[111][85] = 16'h000C;
        rom[111][86] = 16'hFFF9;
        rom[111][87] = 16'h0007;
        rom[111][88] = 16'h0010;
        rom[111][89] = 16'h0013;
        rom[111][90] = 16'hFFFC;
        rom[111][91] = 16'hFFFF;
        rom[111][92] = 16'hFFFE;
        rom[111][93] = 16'hFFF9;
        rom[111][94] = 16'hFFC0;
        rom[111][95] = 16'h000C;
        rom[111][96] = 16'h0016;
        rom[111][97] = 16'h001A;
        rom[111][98] = 16'h000C;
        rom[111][99] = 16'h002B;
        rom[111][100] = 16'h0021;
        rom[111][101] = 16'h0024;
        rom[111][102] = 16'h0016;
        rom[111][103] = 16'h0004;
        rom[111][104] = 16'hFFFD;
        rom[111][105] = 16'hFFF6;
        rom[111][106] = 16'h0014;
        rom[111][107] = 16'h000B;
        rom[111][108] = 16'h0019;
        rom[111][109] = 16'h0011;
        rom[111][110] = 16'h0031;
        rom[111][111] = 16'h0029;
        rom[111][112] = 16'h001B;
        rom[111][113] = 16'hFFF8;
        rom[111][114] = 16'h000E;
        rom[111][115] = 16'hFFFF;
        rom[111][116] = 16'hFFDF;
        rom[111][117] = 16'h000F;
        rom[111][118] = 16'h001C;
        rom[111][119] = 16'h0013;
        rom[111][120] = 16'hFFCB;
        rom[111][121] = 16'h0006;
        rom[111][122] = 16'hFFFC;
        rom[111][123] = 16'hFFBE;
        rom[111][124] = 16'h0009;
        rom[111][125] = 16'h001F;
        rom[111][126] = 16'hFFDD;
        rom[111][127] = 16'hFFE1;
        rom[112][0] = 16'hFFF1;
        rom[112][1] = 16'h0011;
        rom[112][2] = 16'hFFE4;
        rom[112][3] = 16'h0009;
        rom[112][4] = 16'h0016;
        rom[112][5] = 16'hFFCF;
        rom[112][6] = 16'h0012;
        rom[112][7] = 16'hFFDB;
        rom[112][8] = 16'h0010;
        rom[112][9] = 16'h001B;
        rom[112][10] = 16'h0034;
        rom[112][11] = 16'h0029;
        rom[112][12] = 16'h0001;
        rom[112][13] = 16'h000F;
        rom[112][14] = 16'hFFEF;
        rom[112][15] = 16'h0008;
        rom[112][16] = 16'hFFDA;
        rom[112][17] = 16'hFFE1;
        rom[112][18] = 16'hFFCF;
        rom[112][19] = 16'h001D;
        rom[112][20] = 16'h000A;
        rom[112][21] = 16'h000F;
        rom[112][22] = 16'hFFEF;
        rom[112][23] = 16'hFFEA;
        rom[112][24] = 16'h0027;
        rom[112][25] = 16'h0015;
        rom[112][26] = 16'h000E;
        rom[112][27] = 16'h0011;
        rom[112][28] = 16'hFFCA;
        rom[112][29] = 16'hFFBB;
        rom[112][30] = 16'h0029;
        rom[112][31] = 16'hFFFB;
        rom[112][32] = 16'hFFD7;
        rom[112][33] = 16'h003C;
        rom[112][34] = 16'hFFF7;
        rom[112][35] = 16'hFFF3;
        rom[112][36] = 16'hFFF7;
        rom[112][37] = 16'hFFE1;
        rom[112][38] = 16'h000D;
        rom[112][39] = 16'h000F;
        rom[112][40] = 16'hFFEF;
        rom[112][41] = 16'h0021;
        rom[112][42] = 16'hFFD6;
        rom[112][43] = 16'hFFF2;
        rom[112][44] = 16'h001A;
        rom[112][45] = 16'h0001;
        rom[112][46] = 16'hFFE5;
        rom[112][47] = 16'hFFFE;
        rom[112][48] = 16'hFFDC;
        rom[112][49] = 16'hFFB1;
        rom[112][50] = 16'h000E;
        rom[112][51] = 16'hFFF4;
        rom[112][52] = 16'hFFF5;
        rom[112][53] = 16'hFFE2;
        rom[112][54] = 16'h0017;
        rom[112][55] = 16'hFFEE;
        rom[112][56] = 16'hFFF9;
        rom[112][57] = 16'h0011;
        rom[112][58] = 16'hFFFE;
        rom[112][59] = 16'h0013;
        rom[112][60] = 16'h0009;
        rom[112][61] = 16'hFFDA;
        rom[112][62] = 16'h0017;
        rom[112][63] = 16'hFFCD;
        rom[112][64] = 16'hFFD7;
        rom[112][65] = 16'h000C;
        rom[112][66] = 16'hFFF0;
        rom[112][67] = 16'hFFFE;
        rom[112][68] = 16'h0017;
        rom[112][69] = 16'hFFCD;
        rom[112][70] = 16'hFFF4;
        rom[112][71] = 16'hFFE1;
        rom[112][72] = 16'hFFFD;
        rom[112][73] = 16'hFFEF;
        rom[112][74] = 16'h000C;
        rom[112][75] = 16'h0047;
        rom[112][76] = 16'hFFD1;
        rom[112][77] = 16'h001F;
        rom[112][78] = 16'h0035;
        rom[112][79] = 16'h0005;
        rom[112][80] = 16'h0010;
        rom[112][81] = 16'hFFEB;
        rom[112][82] = 16'hFFD3;
        rom[112][83] = 16'h000A;
        rom[112][84] = 16'hFFF9;
        rom[112][85] = 16'h001F;
        rom[112][86] = 16'hFFC7;
        rom[112][87] = 16'h0029;
        rom[112][88] = 16'h0026;
        rom[112][89] = 16'h0027;
        rom[112][90] = 16'hFFC5;
        rom[112][91] = 16'hFFD6;
        rom[112][92] = 16'h0022;
        rom[112][93] = 16'hFFF3;
        rom[112][94] = 16'hFFBD;
        rom[112][95] = 16'hFFF2;
        rom[112][96] = 16'hFFFA;
        rom[112][97] = 16'h0013;
        rom[112][98] = 16'h0006;
        rom[112][99] = 16'h0009;
        rom[112][100] = 16'hFFF6;
        rom[112][101] = 16'hFFC9;
        rom[112][102] = 16'hFFCC;
        rom[112][103] = 16'h001C;
        rom[112][104] = 16'hFFEE;
        rom[112][105] = 16'h000E;
        rom[112][106] = 16'hFFBF;
        rom[112][107] = 16'hFFDC;
        rom[112][108] = 16'hFFE9;
        rom[112][109] = 16'h000F;
        rom[112][110] = 16'hFFD2;
        rom[112][111] = 16'h0006;
        rom[112][112] = 16'h0009;
        rom[112][113] = 16'hFFEC;
        rom[112][114] = 16'h0011;
        rom[112][115] = 16'hFFF0;
        rom[112][116] = 16'h002C;
        rom[112][117] = 16'hFFEC;
        rom[112][118] = 16'hFFFF;
        rom[112][119] = 16'h000C;
        rom[112][120] = 16'h0007;
        rom[112][121] = 16'h001A;
        rom[112][122] = 16'h001C;
        rom[112][123] = 16'hFFE5;
        rom[112][124] = 16'h001E;
        rom[112][125] = 16'h0007;
        rom[112][126] = 16'hFFED;
        rom[112][127] = 16'h001E;
        rom[113][0] = 16'hFFF4;
        rom[113][1] = 16'hFFD9;
        rom[113][2] = 16'h001C;
        rom[113][3] = 16'hFFF2;
        rom[113][4] = 16'h0017;
        rom[113][5] = 16'h0011;
        rom[113][6] = 16'hFFE6;
        rom[113][7] = 16'hFFC3;
        rom[113][8] = 16'hFFD8;
        rom[113][9] = 16'hFFDF;
        rom[113][10] = 16'hFFE9;
        rom[113][11] = 16'h001A;
        rom[113][12] = 16'hFFC5;
        rom[113][13] = 16'h000C;
        rom[113][14] = 16'hFFF2;
        rom[113][15] = 16'h0023;
        rom[113][16] = 16'hFFE1;
        rom[113][17] = 16'h0002;
        rom[113][18] = 16'hFFCF;
        rom[113][19] = 16'hFFFD;
        rom[113][20] = 16'hFFEA;
        rom[113][21] = 16'hFFD1;
        rom[113][22] = 16'hFFF0;
        rom[113][23] = 16'hFFC6;
        rom[113][24] = 16'hFFF9;
        rom[113][25] = 16'h0004;
        rom[113][26] = 16'hFFF3;
        rom[113][27] = 16'hFFFC;
        rom[113][28] = 16'hFFF2;
        rom[113][29] = 16'hFFEC;
        rom[113][30] = 16'hFFE8;
        rom[113][31] = 16'hFFC2;
        rom[113][32] = 16'h0015;
        rom[113][33] = 16'hFFD5;
        rom[113][34] = 16'hFFF9;
        rom[113][35] = 16'h0028;
        rom[113][36] = 16'hFFA0;
        rom[113][37] = 16'hFFFE;
        rom[113][38] = 16'hFFF0;
        rom[113][39] = 16'hFFFF;
        rom[113][40] = 16'hFFEC;
        rom[113][41] = 16'hFFF6;
        rom[113][42] = 16'hFFD1;
        rom[113][43] = 16'h0006;
        rom[113][44] = 16'h001C;
        rom[113][45] = 16'h0017;
        rom[113][46] = 16'hFFE2;
        rom[113][47] = 16'hFFDD;
        rom[113][48] = 16'h0004;
        rom[113][49] = 16'h000A;
        rom[113][50] = 16'h0019;
        rom[113][51] = 16'h0005;
        rom[113][52] = 16'h0009;
        rom[113][53] = 16'h0027;
        rom[113][54] = 16'h0007;
        rom[113][55] = 16'hFFF9;
        rom[113][56] = 16'hFFF3;
        rom[113][57] = 16'h0033;
        rom[113][58] = 16'hFFCB;
        rom[113][59] = 16'hFFF9;
        rom[113][60] = 16'h000E;
        rom[113][61] = 16'hFFF2;
        rom[113][62] = 16'h0008;
        rom[113][63] = 16'hFFE1;
        rom[113][64] = 16'h0017;
        rom[113][65] = 16'hFFCD;
        rom[113][66] = 16'h001F;
        rom[113][67] = 16'h0002;
        rom[113][68] = 16'h002C;
        rom[113][69] = 16'hFFD8;
        rom[113][70] = 16'h000A;
        rom[113][71] = 16'h0014;
        rom[113][72] = 16'hFFF9;
        rom[113][73] = 16'h000D;
        rom[113][74] = 16'hFFB8;
        rom[113][75] = 16'hFFC6;
        rom[113][76] = 16'hFFF9;
        rom[113][77] = 16'hFFF7;
        rom[113][78] = 16'h0001;
        rom[113][79] = 16'hFFD5;
        rom[113][80] = 16'hFFDD;
        rom[113][81] = 16'hFFFA;
        rom[113][82] = 16'h000C;
        rom[113][83] = 16'hFFE5;
        rom[113][84] = 16'h0006;
        rom[113][85] = 16'h0006;
        rom[113][86] = 16'h0016;
        rom[113][87] = 16'hFFEA;
        rom[113][88] = 16'hFFF7;
        rom[113][89] = 16'h001A;
        rom[113][90] = 16'hFFFE;
        rom[113][91] = 16'hFFD7;
        rom[113][92] = 16'hFFEF;
        rom[113][93] = 16'hFFD9;
        rom[113][94] = 16'hFFC8;
        rom[113][95] = 16'hFFCD;
        rom[113][96] = 16'h0013;
        rom[113][97] = 16'hFFE5;
        rom[113][98] = 16'h0000;
        rom[113][99] = 16'hFFBF;
        rom[113][100] = 16'hFFD8;
        rom[113][101] = 16'hFFEA;
        rom[113][102] = 16'hFFC7;
        rom[113][103] = 16'hFFCD;
        rom[113][104] = 16'h0025;
        rom[113][105] = 16'h0005;
        rom[113][106] = 16'hFFFB;
        rom[113][107] = 16'h001D;
        rom[113][108] = 16'h0000;
        rom[113][109] = 16'hFFEC;
        rom[113][110] = 16'h0024;
        rom[113][111] = 16'hFFF3;
        rom[113][112] = 16'hFFEF;
        rom[113][113] = 16'hFFC4;
        rom[113][114] = 16'h0008;
        rom[113][115] = 16'hFFE2;
        rom[113][116] = 16'hFFB4;
        rom[113][117] = 16'hFFE5;
        rom[113][118] = 16'hFFFE;
        rom[113][119] = 16'h000C;
        rom[113][120] = 16'h0032;
        rom[113][121] = 16'hFFF2;
        rom[113][122] = 16'h0009;
        rom[113][123] = 16'h0011;
        rom[113][124] = 16'h0016;
        rom[113][125] = 16'hFFEF;
        rom[113][126] = 16'hFFF8;
        rom[113][127] = 16'hFFFA;
        rom[114][0] = 16'hFFE6;
        rom[114][1] = 16'hFFF8;
        rom[114][2] = 16'hFFB8;
        rom[114][3] = 16'h0012;
        rom[114][4] = 16'h0002;
        rom[114][5] = 16'hFFFF;
        rom[114][6] = 16'hFFFB;
        rom[114][7] = 16'hFFE8;
        rom[114][8] = 16'hFFF5;
        rom[114][9] = 16'hFFCA;
        rom[114][10] = 16'hFFDA;
        rom[114][11] = 16'h0024;
        rom[114][12] = 16'h000D;
        rom[114][13] = 16'hFFE1;
        rom[114][14] = 16'hFFC3;
        rom[114][15] = 16'h002A;
        rom[114][16] = 16'hFFFF;
        rom[114][17] = 16'hFFD4;
        rom[114][18] = 16'h0011;
        rom[114][19] = 16'hFFFF;
        rom[114][20] = 16'hFFD4;
        rom[114][21] = 16'h0011;
        rom[114][22] = 16'h000A;
        rom[114][23] = 16'hFFC4;
        rom[114][24] = 16'h001B;
        rom[114][25] = 16'hFFDA;
        rom[114][26] = 16'hFFFB;
        rom[114][27] = 16'hFFF6;
        rom[114][28] = 16'h0010;
        rom[114][29] = 16'hFFFF;
        rom[114][30] = 16'h0016;
        rom[114][31] = 16'hFFFB;
        rom[114][32] = 16'hFFD2;
        rom[114][33] = 16'h000E;
        rom[114][34] = 16'hFFE1;
        rom[114][35] = 16'h0020;
        rom[114][36] = 16'h000B;
        rom[114][37] = 16'h000B;
        rom[114][38] = 16'hFFA7;
        rom[114][39] = 16'h000C;
        rom[114][40] = 16'hFFB8;
        rom[114][41] = 16'hFFE3;
        rom[114][42] = 16'h0029;
        rom[114][43] = 16'h0022;
        rom[114][44] = 16'h0012;
        rom[114][45] = 16'hFFE9;
        rom[114][46] = 16'h0003;
        rom[114][47] = 16'hFFFE;
        rom[114][48] = 16'hFFB9;
        rom[114][49] = 16'hFFD7;
        rom[114][50] = 16'hFFD1;
        rom[114][51] = 16'hFFD1;
        rom[114][52] = 16'h0001;
        rom[114][53] = 16'h0002;
        rom[114][54] = 16'h000C;
        rom[114][55] = 16'h000D;
        rom[114][56] = 16'hFFF4;
        rom[114][57] = 16'hFFCE;
        rom[114][58] = 16'h0021;
        rom[114][59] = 16'h0002;
        rom[114][60] = 16'h001B;
        rom[114][61] = 16'hFFFB;
        rom[114][62] = 16'h0010;
        rom[114][63] = 16'hFFDD;
        rom[114][64] = 16'h0022;
        rom[114][65] = 16'h0016;
        rom[114][66] = 16'h0019;
        rom[114][67] = 16'hFFEF;
        rom[114][68] = 16'hFFF1;
        rom[114][69] = 16'h0007;
        rom[114][70] = 16'hFFC5;
        rom[114][71] = 16'h0013;
        rom[114][72] = 16'hFFEE;
        rom[114][73] = 16'hFFE5;
        rom[114][74] = 16'hFFE8;
        rom[114][75] = 16'hFFF7;
        rom[114][76] = 16'h0032;
        rom[114][77] = 16'h0018;
        rom[114][78] = 16'h0008;
        rom[114][79] = 16'h0024;
        rom[114][80] = 16'hFFEF;
        rom[114][81] = 16'h001E;
        rom[114][82] = 16'hFFD4;
        rom[114][83] = 16'h0031;
        rom[114][84] = 16'h0002;
        rom[114][85] = 16'h001A;
        rom[114][86] = 16'hFFDF;
        rom[114][87] = 16'h0005;
        rom[114][88] = 16'hFF9A;
        rom[114][89] = 16'h000A;
        rom[114][90] = 16'hFFC1;
        rom[114][91] = 16'h0013;
        rom[114][92] = 16'h0007;
        rom[114][93] = 16'h0002;
        rom[114][94] = 16'hFFED;
        rom[114][95] = 16'h000A;
        rom[114][96] = 16'hFFF5;
        rom[114][97] = 16'hFFAC;
        rom[114][98] = 16'h0004;
        rom[114][99] = 16'h0015;
        rom[114][100] = 16'h0016;
        rom[114][101] = 16'hFFF1;
        rom[114][102] = 16'hFFD8;
        rom[114][103] = 16'hFFF3;
        rom[114][104] = 16'h0015;
        rom[114][105] = 16'hFFD3;
        rom[114][106] = 16'hFFED;
        rom[114][107] = 16'h001A;
        rom[114][108] = 16'hFFD8;
        rom[114][109] = 16'h001B;
        rom[114][110] = 16'h0014;
        rom[114][111] = 16'h002E;
        rom[114][112] = 16'hFFFF;
        rom[114][113] = 16'h0011;
        rom[114][114] = 16'hFFF0;
        rom[114][115] = 16'hFFF4;
        rom[114][116] = 16'hFFF9;
        rom[114][117] = 16'hFFEA;
        rom[114][118] = 16'h0013;
        rom[114][119] = 16'hFFF2;
        rom[114][120] = 16'h0002;
        rom[114][121] = 16'hFFE3;
        rom[114][122] = 16'h0024;
        rom[114][123] = 16'hFFE5;
        rom[114][124] = 16'h0025;
        rom[114][125] = 16'h0028;
        rom[114][126] = 16'hFFE4;
        rom[114][127] = 16'h0003;
        rom[115][0] = 16'h0000;
        rom[115][1] = 16'h0001;
        rom[115][2] = 16'hFFC4;
        rom[115][3] = 16'hFFF5;
        rom[115][4] = 16'hFFED;
        rom[115][5] = 16'hFFC0;
        rom[115][6] = 16'hFFF4;
        rom[115][7] = 16'h0013;
        rom[115][8] = 16'h0039;
        rom[115][9] = 16'hFFF4;
        rom[115][10] = 16'h003C;
        rom[115][11] = 16'h000B;
        rom[115][12] = 16'h0007;
        rom[115][13] = 16'h0015;
        rom[115][14] = 16'hFFB0;
        rom[115][15] = 16'hFFD2;
        rom[115][16] = 16'h001A;
        rom[115][17] = 16'h0023;
        rom[115][18] = 16'hFFB8;
        rom[115][19] = 16'h0017;
        rom[115][20] = 16'h0045;
        rom[115][21] = 16'h0004;
        rom[115][22] = 16'hFFE5;
        rom[115][23] = 16'h000C;
        rom[115][24] = 16'h0009;
        rom[115][25] = 16'hFFD0;
        rom[115][26] = 16'h0000;
        rom[115][27] = 16'h0006;
        rom[115][28] = 16'hFFF2;
        rom[115][29] = 16'hFFDA;
        rom[115][30] = 16'hFFDA;
        rom[115][31] = 16'h003D;
        rom[115][32] = 16'hFFD3;
        rom[115][33] = 16'h0029;
        rom[115][34] = 16'h0003;
        rom[115][35] = 16'hFFC8;
        rom[115][36] = 16'h0006;
        rom[115][37] = 16'hFFEA;
        rom[115][38] = 16'hFFD7;
        rom[115][39] = 16'hFFF9;
        rom[115][40] = 16'hFFEA;
        rom[115][41] = 16'h0003;
        rom[115][42] = 16'hFFFB;
        rom[115][43] = 16'hFFE4;
        rom[115][44] = 16'h0018;
        rom[115][45] = 16'hFFB7;
        rom[115][46] = 16'h000B;
        rom[115][47] = 16'h001F;
        rom[115][48] = 16'hFFD4;
        rom[115][49] = 16'hFFF6;
        rom[115][50] = 16'hFFF1;
        rom[115][51] = 16'h0002;
        rom[115][52] = 16'hFFEA;
        rom[115][53] = 16'hFFD2;
        rom[115][54] = 16'hFFEF;
        rom[115][55] = 16'hFFD3;
        rom[115][56] = 16'hFFED;
        rom[115][57] = 16'hFFE8;
        rom[115][58] = 16'h0021;
        rom[115][59] = 16'h0004;
        rom[115][60] = 16'hFFF9;
        rom[115][61] = 16'h0009;
        rom[115][62] = 16'h000C;
        rom[115][63] = 16'hFFAA;
        rom[115][64] = 16'h0029;
        rom[115][65] = 16'h0008;
        rom[115][66] = 16'hFFEE;
        rom[115][67] = 16'hFFED;
        rom[115][68] = 16'hFFEA;
        rom[115][69] = 16'hFFF8;
        rom[115][70] = 16'hFFED;
        rom[115][71] = 16'hFFF9;
        rom[115][72] = 16'hFFFF;
        rom[115][73] = 16'hFFE5;
        rom[115][74] = 16'h0022;
        rom[115][75] = 16'h0007;
        rom[115][76] = 16'h000C;
        rom[115][77] = 16'h0011;
        rom[115][78] = 16'h0024;
        rom[115][79] = 16'h0014;
        rom[115][80] = 16'hFFED;
        rom[115][81] = 16'h0016;
        rom[115][82] = 16'h001E;
        rom[115][83] = 16'h0026;
        rom[115][84] = 16'hFFE8;
        rom[115][85] = 16'hFFE8;
        rom[115][86] = 16'hFFCB;
        rom[115][87] = 16'h000F;
        rom[115][88] = 16'h0018;
        rom[115][89] = 16'hFFDA;
        rom[115][90] = 16'hFFFC;
        rom[115][91] = 16'hFFEA;
        rom[115][92] = 16'h002C;
        rom[115][93] = 16'hFFDD;
        rom[115][94] = 16'h000B;
        rom[115][95] = 16'hFFEC;
        rom[115][96] = 16'hFFE8;
        rom[115][97] = 16'hFFE9;
        rom[115][98] = 16'h0042;
        rom[115][99] = 16'h000C;
        rom[115][100] = 16'h0008;
        rom[115][101] = 16'h0047;
        rom[115][102] = 16'hFFF6;
        rom[115][103] = 16'hFFF9;
        rom[115][104] = 16'h0002;
        rom[115][105] = 16'hFFDF;
        rom[115][106] = 16'hFFFA;
        rom[115][107] = 16'hFFC7;
        rom[115][108] = 16'hFFE6;
        rom[115][109] = 16'h0001;
        rom[115][110] = 16'hFFD2;
        rom[115][111] = 16'hFFF8;
        rom[115][112] = 16'h0015;
        rom[115][113] = 16'hFFB2;
        rom[115][114] = 16'hFFEF;
        rom[115][115] = 16'h0011;
        rom[115][116] = 16'hFFFE;
        rom[115][117] = 16'hFFDF;
        rom[115][118] = 16'hFFDC;
        rom[115][119] = 16'h0000;
        rom[115][120] = 16'h0000;
        rom[115][121] = 16'hFFDE;
        rom[115][122] = 16'h000E;
        rom[115][123] = 16'hFFFE;
        rom[115][124] = 16'hFFF8;
        rom[115][125] = 16'h001B;
        rom[115][126] = 16'hFFD2;
        rom[115][127] = 16'hFFB1;
        rom[116][0] = 16'hFFF4;
        rom[116][1] = 16'hFFF9;
        rom[116][2] = 16'h0023;
        rom[116][3] = 16'h0016;
        rom[116][4] = 16'h0005;
        rom[116][5] = 16'hFFFE;
        rom[116][6] = 16'hFFEF;
        rom[116][7] = 16'hFFF6;
        rom[116][8] = 16'hFFC3;
        rom[116][9] = 16'h0003;
        rom[116][10] = 16'h0011;
        rom[116][11] = 16'h0036;
        rom[116][12] = 16'h0006;
        rom[116][13] = 16'h0019;
        rom[116][14] = 16'h0026;
        rom[116][15] = 16'h0025;
        rom[116][16] = 16'hFFFA;
        rom[116][17] = 16'hFFD2;
        rom[116][18] = 16'hFFDA;
        rom[116][19] = 16'hFFF4;
        rom[116][20] = 16'h0020;
        rom[116][21] = 16'hFFD2;
        rom[116][22] = 16'h0003;
        rom[116][23] = 16'hFFF4;
        rom[116][24] = 16'hFFED;
        rom[116][25] = 16'h0003;
        rom[116][26] = 16'h000B;
        rom[116][27] = 16'h0011;
        rom[116][28] = 16'h0007;
        rom[116][29] = 16'h0020;
        rom[116][30] = 16'hFFCF;
        rom[116][31] = 16'hFFAD;
        rom[116][32] = 16'h001E;
        rom[116][33] = 16'hFFD9;
        rom[116][34] = 16'hFFC6;
        rom[116][35] = 16'h0016;
        rom[116][36] = 16'hFFED;
        rom[116][37] = 16'hFFF9;
        rom[116][38] = 16'h0000;
        rom[116][39] = 16'hFFC4;
        rom[116][40] = 16'hFFF0;
        rom[116][41] = 16'hFFFF;
        rom[116][42] = 16'hFFEF;
        rom[116][43] = 16'hFFED;
        rom[116][44] = 16'hFFD9;
        rom[116][45] = 16'h000B;
        rom[116][46] = 16'hFFEF;
        rom[116][47] = 16'hFFDC;
        rom[116][48] = 16'h0013;
        rom[116][49] = 16'hFFF2;
        rom[116][50] = 16'h002A;
        rom[116][51] = 16'hFFC8;
        rom[116][52] = 16'hFFDB;
        rom[116][53] = 16'h0001;
        rom[116][54] = 16'h0009;
        rom[116][55] = 16'hFFE2;
        rom[116][56] = 16'h0012;
        rom[116][57] = 16'h001F;
        rom[116][58] = 16'hFFC9;
        rom[116][59] = 16'hFFFC;
        rom[116][60] = 16'hFFF9;
        rom[116][61] = 16'h001B;
        rom[116][62] = 16'hFFE9;
        rom[116][63] = 16'hFFF4;
        rom[116][64] = 16'hFFD4;
        rom[116][65] = 16'hFFD7;
        rom[116][66] = 16'h0016;
        rom[116][67] = 16'h0013;
        rom[116][68] = 16'h000B;
        rom[116][69] = 16'h0007;
        rom[116][70] = 16'h0034;
        rom[116][71] = 16'hFFF1;
        rom[116][72] = 16'h000C;
        rom[116][73] = 16'h0018;
        rom[116][74] = 16'hFFB0;
        rom[116][75] = 16'hFFD6;
        rom[116][76] = 16'hFFFD;
        rom[116][77] = 16'hFFE5;
        rom[116][78] = 16'h0023;
        rom[116][79] = 16'hFFB0;
        rom[116][80] = 16'h0004;
        rom[116][81] = 16'h0023;
        rom[116][82] = 16'h0007;
        rom[116][83] = 16'h0016;
        rom[116][84] = 16'h0010;
        rom[116][85] = 16'hFFE7;
        rom[116][86] = 16'hFFF4;
        rom[116][87] = 16'hFFE9;
        rom[116][88] = 16'h0004;
        rom[116][89] = 16'h001A;
        rom[116][90] = 16'h0009;
        rom[116][91] = 16'hFFDD;
        rom[116][92] = 16'hFFD2;
        rom[116][93] = 16'h0032;
        rom[116][94] = 16'hFFD6;
        rom[116][95] = 16'hFFF9;
        rom[116][96] = 16'h002D;
        rom[116][97] = 16'h000C;
        rom[116][98] = 16'hFFE4;
        rom[116][99] = 16'hFFF4;
        rom[116][100] = 16'hFFE6;
        rom[116][101] = 16'hFFEF;
        rom[116][102] = 16'h000E;
        rom[116][103] = 16'h0004;
        rom[116][104] = 16'h0007;
        rom[116][105] = 16'hFFC1;
        rom[116][106] = 16'hFFED;
        rom[116][107] = 16'h001C;
        rom[116][108] = 16'hFFDE;
        rom[116][109] = 16'h0024;
        rom[116][110] = 16'h0014;
        rom[116][111] = 16'h002B;
        rom[116][112] = 16'h002B;
        rom[116][113] = 16'hFFEA;
        rom[116][114] = 16'h000C;
        rom[116][115] = 16'hFFEF;
        rom[116][116] = 16'hFFBA;
        rom[116][117] = 16'hFFE8;
        rom[116][118] = 16'hFFD7;
        rom[116][119] = 16'h001F;
        rom[116][120] = 16'hFFE5;
        rom[116][121] = 16'hFFE8;
        rom[116][122] = 16'h001A;
        rom[116][123] = 16'hFFBE;
        rom[116][124] = 16'h000E;
        rom[116][125] = 16'hFFF5;
        rom[116][126] = 16'h000B;
        rom[116][127] = 16'h0001;
        rom[117][0] = 16'h0023;
        rom[117][1] = 16'hFFDF;
        rom[117][2] = 16'h0000;
        rom[117][3] = 16'h0028;
        rom[117][4] = 16'hFFE9;
        rom[117][5] = 16'hFFEA;
        rom[117][6] = 16'hFFEE;
        rom[117][7] = 16'h0012;
        rom[117][8] = 16'hFFD3;
        rom[117][9] = 16'h000F;
        rom[117][10] = 16'hFFF1;
        rom[117][11] = 16'hFFEC;
        rom[117][12] = 16'hFFCB;
        rom[117][13] = 16'hFFEA;
        rom[117][14] = 16'hFFDC;
        rom[117][15] = 16'h0009;
        rom[117][16] = 16'hFFFB;
        rom[117][17] = 16'h0004;
        rom[117][18] = 16'h0011;
        rom[117][19] = 16'hFFC9;
        rom[117][20] = 16'h0004;
        rom[117][21] = 16'h0005;
        rom[117][22] = 16'hFFEA;
        rom[117][23] = 16'h0026;
        rom[117][24] = 16'h000F;
        rom[117][25] = 16'h0009;
        rom[117][26] = 16'hFFDB;
        rom[117][27] = 16'hFFCC;
        rom[117][28] = 16'hFFF5;
        rom[117][29] = 16'hFFD7;
        rom[117][30] = 16'hFFFF;
        rom[117][31] = 16'h001A;
        rom[117][32] = 16'h0006;
        rom[117][33] = 16'hFFFC;
        rom[117][34] = 16'h0010;
        rom[117][35] = 16'h0007;
        rom[117][36] = 16'h0023;
        rom[117][37] = 16'hFFCE;
        rom[117][38] = 16'h0033;
        rom[117][39] = 16'hFFEF;
        rom[117][40] = 16'hFFF9;
        rom[117][41] = 16'h001E;
        rom[117][42] = 16'hFFE2;
        rom[117][43] = 16'h0017;
        rom[117][44] = 16'h001C;
        rom[117][45] = 16'hFFFA;
        rom[117][46] = 16'h0033;
        rom[117][47] = 16'hFFF9;
        rom[117][48] = 16'h000B;
        rom[117][49] = 16'hFFF9;
        rom[117][50] = 16'h0012;
        rom[117][51] = 16'h000A;
        rom[117][52] = 16'hFFDC;
        rom[117][53] = 16'h0002;
        rom[117][54] = 16'hFFC7;
        rom[117][55] = 16'h0007;
        rom[117][56] = 16'hFFD0;
        rom[117][57] = 16'h0003;
        rom[117][58] = 16'hFFE2;
        rom[117][59] = 16'h0003;
        rom[117][60] = 16'hFFEB;
        rom[117][61] = 16'hFFFC;
        rom[117][62] = 16'hFFEF;
        rom[117][63] = 16'h000E;
        rom[117][64] = 16'h0024;
        rom[117][65] = 16'h0016;
        rom[117][66] = 16'hFFE1;
        rom[117][67] = 16'hFFBF;
        rom[117][68] = 16'h0010;
        rom[117][69] = 16'hFFCF;
        rom[117][70] = 16'h0002;
        rom[117][71] = 16'hFFD7;
        rom[117][72] = 16'h0012;
        rom[117][73] = 16'hFFF4;
        rom[117][74] = 16'h001B;
        rom[117][75] = 16'h0003;
        rom[117][76] = 16'h0009;
        rom[117][77] = 16'hFFC3;
        rom[117][78] = 16'hFFE3;
        rom[117][79] = 16'hFFD5;
        rom[117][80] = 16'h0003;
        rom[117][81] = 16'hFFBF;
        rom[117][82] = 16'h0007;
        rom[117][83] = 16'hFFDF;
        rom[117][84] = 16'hFFFF;
        rom[117][85] = 16'h0016;
        rom[117][86] = 16'h0017;
        rom[117][87] = 16'h0009;
        rom[117][88] = 16'h0033;
        rom[117][89] = 16'hFFD4;
        rom[117][90] = 16'hFFFD;
        rom[117][91] = 16'hFFE6;
        rom[117][92] = 16'hFFFA;
        rom[117][93] = 16'hFFF2;
        rom[117][94] = 16'hFFF8;
        rom[117][95] = 16'hFFCD;
        rom[117][96] = 16'h0000;
        rom[117][97] = 16'hFFF4;
        rom[117][98] = 16'hFFF1;
        rom[117][99] = 16'hFFE1;
        rom[117][100] = 16'hFFDA;
        rom[117][101] = 16'h002C;
        rom[117][102] = 16'hFFD4;
        rom[117][103] = 16'hFFDD;
        rom[117][104] = 16'h0007;
        rom[117][105] = 16'hFFCE;
        rom[117][106] = 16'h0012;
        rom[117][107] = 16'hFFEB;
        rom[117][108] = 16'hFFCD;
        rom[117][109] = 16'hFFF6;
        rom[117][110] = 16'h0022;
        rom[117][111] = 16'hFFB2;
        rom[117][112] = 16'hFFFD;
        rom[117][113] = 16'hFFC4;
        rom[117][114] = 16'hFFD6;
        rom[117][115] = 16'h001A;
        rom[117][116] = 16'h001F;
        rom[117][117] = 16'hFFF2;
        rom[117][118] = 16'h0027;
        rom[117][119] = 16'h0012;
        rom[117][120] = 16'h0010;
        rom[117][121] = 16'h0001;
        rom[117][122] = 16'hFFF4;
        rom[117][123] = 16'h0037;
        rom[117][124] = 16'hFFCD;
        rom[117][125] = 16'h0011;
        rom[117][126] = 16'hFFC3;
        rom[117][127] = 16'hFFC3;
        rom[118][0] = 16'h001F;
        rom[118][1] = 16'h0011;
        rom[118][2] = 16'hFFEF;
        rom[118][3] = 16'h002E;
        rom[118][4] = 16'h0013;
        rom[118][5] = 16'hFFFE;
        rom[118][6] = 16'hFFCD;
        rom[118][7] = 16'h0022;
        rom[118][8] = 16'h0009;
        rom[118][9] = 16'h002E;
        rom[118][10] = 16'h0014;
        rom[118][11] = 16'h0016;
        rom[118][12] = 16'hFFE4;
        rom[118][13] = 16'hFFEF;
        rom[118][14] = 16'h0009;
        rom[118][15] = 16'hFFE5;
        rom[118][16] = 16'hFFAC;
        rom[118][17] = 16'hFFF6;
        rom[118][18] = 16'h002C;
        rom[118][19] = 16'hFFF8;
        rom[118][20] = 16'h0029;
        rom[118][21] = 16'h000D;
        rom[118][22] = 16'hFFF8;
        rom[118][23] = 16'h0027;
        rom[118][24] = 16'hFFFE;
        rom[118][25] = 16'h002C;
        rom[118][26] = 16'hFFF1;
        rom[118][27] = 16'hFFE8;
        rom[118][28] = 16'h0018;
        rom[118][29] = 16'hFFE5;
        rom[118][30] = 16'hFFE6;
        rom[118][31] = 16'hFFEA;
        rom[118][32] = 16'hFFEF;
        rom[118][33] = 16'h001A;
        rom[118][34] = 16'hFFDC;
        rom[118][35] = 16'hFFFF;
        rom[118][36] = 16'hFFF5;
        rom[118][37] = 16'hFFEF;
        rom[118][38] = 16'h0028;
        rom[118][39] = 16'hFFF4;
        rom[118][40] = 16'hFFF8;
        rom[118][41] = 16'hFFEA;
        rom[118][42] = 16'h0018;
        rom[118][43] = 16'hFFD2;
        rom[118][44] = 16'hFFC0;
        rom[118][45] = 16'h0007;
        rom[118][46] = 16'hFFEF;
        rom[118][47] = 16'hFFE1;
        rom[118][48] = 16'hFFD5;
        rom[118][49] = 16'h0008;
        rom[118][50] = 16'h0003;
        rom[118][51] = 16'hFFF4;
        rom[118][52] = 16'h0014;
        rom[118][53] = 16'hFFF4;
        rom[118][54] = 16'hFFFF;
        rom[118][55] = 16'h001B;
        rom[118][56] = 16'hFFFC;
        rom[118][57] = 16'hFFFE;
        rom[118][58] = 16'hFFD7;
        rom[118][59] = 16'h0016;
        rom[118][60] = 16'hFFBD;
        rom[118][61] = 16'hFFBC;
        rom[118][62] = 16'h0006;
        rom[118][63] = 16'hFFDA;
        rom[118][64] = 16'hFFEA;
        rom[118][65] = 16'hFFE6;
        rom[118][66] = 16'h002E;
        rom[118][67] = 16'h0012;
        rom[118][68] = 16'hFFFC;
        rom[118][69] = 16'h0019;
        rom[118][70] = 16'hFFF7;
        rom[118][71] = 16'h0008;
        rom[118][72] = 16'hFFF6;
        rom[118][73] = 16'h0008;
        rom[118][74] = 16'h0003;
        rom[118][75] = 16'h0032;
        rom[118][76] = 16'h0012;
        rom[118][77] = 16'h0006;
        rom[118][78] = 16'hFFF2;
        rom[118][79] = 16'hFFD2;
        rom[118][80] = 16'h0013;
        rom[118][81] = 16'hFFF0;
        rom[118][82] = 16'h001F;
        rom[118][83] = 16'hFFF8;
        rom[118][84] = 16'hFFCA;
        rom[118][85] = 16'hFFF2;
        rom[118][86] = 16'h0010;
        rom[118][87] = 16'h0012;
        rom[118][88] = 16'h003C;
        rom[118][89] = 16'hFFFD;
        rom[118][90] = 16'h0013;
        rom[118][91] = 16'hFFF9;
        rom[118][92] = 16'hFFFB;
        rom[118][93] = 16'h0011;
        rom[118][94] = 16'h0002;
        rom[118][95] = 16'h000D;
        rom[118][96] = 16'h002B;
        rom[118][97] = 16'hFFFA;
        rom[118][98] = 16'hFFC8;
        rom[118][99] = 16'hFFB5;
        rom[118][100] = 16'h0005;
        rom[118][101] = 16'h0026;
        rom[118][102] = 16'h000E;
        rom[118][103] = 16'h0016;
        rom[118][104] = 16'h000F;
        rom[118][105] = 16'hFFE4;
        rom[118][106] = 16'hFFF1;
        rom[118][107] = 16'h0024;
        rom[118][108] = 16'hFFAD;
        rom[118][109] = 16'hFFED;
        rom[118][110] = 16'hFFF0;
        rom[118][111] = 16'h0017;
        rom[118][112] = 16'h0001;
        rom[118][113] = 16'hFFEE;
        rom[118][114] = 16'hFFD1;
        rom[118][115] = 16'hFFCF;
        rom[118][116] = 16'h0002;
        rom[118][117] = 16'h0000;
        rom[118][118] = 16'h0007;
        rom[118][119] = 16'h001B;
        rom[118][120] = 16'hFFE3;
        rom[118][121] = 16'h001C;
        rom[118][122] = 16'hFFFE;
        rom[118][123] = 16'hFFE1;
        rom[118][124] = 16'h0007;
        rom[118][125] = 16'h0029;
        rom[118][126] = 16'hFFFB;
        rom[118][127] = 16'h0010;
        rom[119][0] = 16'hFFDC;
        rom[119][1] = 16'h0025;
        rom[119][2] = 16'hFFF2;
        rom[119][3] = 16'hFFDC;
        rom[119][4] = 16'h0034;
        rom[119][5] = 16'h001D;
        rom[119][6] = 16'h001D;
        rom[119][7] = 16'h0017;
        rom[119][8] = 16'h000A;
        rom[119][9] = 16'hFFD2;
        rom[119][10] = 16'hFFFB;
        rom[119][11] = 16'hFFD2;
        rom[119][12] = 16'hFFEF;
        rom[119][13] = 16'hFFE5;
        rom[119][14] = 16'hFFF5;
        rom[119][15] = 16'h0000;
        rom[119][16] = 16'h0023;
        rom[119][17] = 16'hFFD8;
        rom[119][18] = 16'hFFFF;
        rom[119][19] = 16'hFFEC;
        rom[119][20] = 16'hFFEA;
        rom[119][21] = 16'hFFEA;
        rom[119][22] = 16'h000B;
        rom[119][23] = 16'hFFFE;
        rom[119][24] = 16'hFFE8;
        rom[119][25] = 16'h0012;
        rom[119][26] = 16'hFFEE;
        rom[119][27] = 16'h001F;
        rom[119][28] = 16'h0010;
        rom[119][29] = 16'hFFF8;
        rom[119][30] = 16'hFFFE;
        rom[119][31] = 16'hFFFE;
        rom[119][32] = 16'h0018;
        rom[119][33] = 16'hFFDA;
        rom[119][34] = 16'hFFE7;
        rom[119][35] = 16'h0003;
        rom[119][36] = 16'h0012;
        rom[119][37] = 16'hFFEC;
        rom[119][38] = 16'hFFEC;
        rom[119][39] = 16'h0002;
        rom[119][40] = 16'h0029;
        rom[119][41] = 16'h000C;
        rom[119][42] = 16'hFFB8;
        rom[119][43] = 16'hFFFE;
        rom[119][44] = 16'hFFFD;
        rom[119][45] = 16'hFFF9;
        rom[119][46] = 16'h000F;
        rom[119][47] = 16'h0002;
        rom[119][48] = 16'h0020;
        rom[119][49] = 16'h0013;
        rom[119][50] = 16'hFFF9;
        rom[119][51] = 16'h0001;
        rom[119][52] = 16'h000C;
        rom[119][53] = 16'hFFF9;
        rom[119][54] = 16'h001E;
        rom[119][55] = 16'h001C;
        rom[119][56] = 16'hFFF0;
        rom[119][57] = 16'hFFFF;
        rom[119][58] = 16'hFFDC;
        rom[119][59] = 16'hFFE6;
        rom[119][60] = 16'hFFF2;
        rom[119][61] = 16'hFFDC;
        rom[119][62] = 16'h002C;
        rom[119][63] = 16'h001A;
        rom[119][64] = 16'hFFF2;
        rom[119][65] = 16'h0038;
        rom[119][66] = 16'h0047;
        rom[119][67] = 16'hFFFF;
        rom[119][68] = 16'h000A;
        rom[119][69] = 16'h0002;
        rom[119][70] = 16'h0002;
        rom[119][71] = 16'h0027;
        rom[119][72] = 16'hFFE0;
        rom[119][73] = 16'h001F;
        rom[119][74] = 16'h0016;
        rom[119][75] = 16'hFFEB;
        rom[119][76] = 16'hFFD5;
        rom[119][77] = 16'hFFF9;
        rom[119][78] = 16'h001C;
        rom[119][79] = 16'h003F;
        rom[119][80] = 16'h0001;
        rom[119][81] = 16'h0002;
        rom[119][82] = 16'h0006;
        rom[119][83] = 16'h0014;
        rom[119][84] = 16'h002C;
        rom[119][85] = 16'h0015;
        rom[119][86] = 16'hFFFA;
        rom[119][87] = 16'h0011;
        rom[119][88] = 16'hFFFC;
        rom[119][89] = 16'h001B;
        rom[119][90] = 16'h000F;
        rom[119][91] = 16'h000A;
        rom[119][92] = 16'hFFB3;
        rom[119][93] = 16'hFFE1;
        rom[119][94] = 16'hFFCD;
        rom[119][95] = 16'h0010;
        rom[119][96] = 16'h001C;
        rom[119][97] = 16'h002A;
        rom[119][98] = 16'hFFFE;
        rom[119][99] = 16'h0011;
        rom[119][100] = 16'h001D;
        rom[119][101] = 16'h0017;
        rom[119][102] = 16'h0010;
        rom[119][103] = 16'hFFF8;
        rom[119][104] = 16'h000A;
        rom[119][105] = 16'hFFD5;
        rom[119][106] = 16'h0002;
        rom[119][107] = 16'h000A;
        rom[119][108] = 16'h0002;
        rom[119][109] = 16'hFFEC;
        rom[119][110] = 16'h0028;
        rom[119][111] = 16'h000C;
        rom[119][112] = 16'h0002;
        rom[119][113] = 16'h0007;
        rom[119][114] = 16'h0001;
        rom[119][115] = 16'h0024;
        rom[119][116] = 16'hFFDC;
        rom[119][117] = 16'h000B;
        rom[119][118] = 16'h0037;
        rom[119][119] = 16'h001D;
        rom[119][120] = 16'hFFE4;
        rom[119][121] = 16'hFFDF;
        rom[119][122] = 16'hFF9C;
        rom[119][123] = 16'hFFBD;
        rom[119][124] = 16'h0037;
        rom[119][125] = 16'h0028;
        rom[119][126] = 16'hFFF6;
        rom[119][127] = 16'hFFCE;
        rom[120][0] = 16'h0002;
        rom[120][1] = 16'hFFE4;
        rom[120][2] = 16'h0002;
        rom[120][3] = 16'hFFD4;
        rom[120][4] = 16'hFFFC;
        rom[120][5] = 16'hFFE9;
        rom[120][6] = 16'hFFEA;
        rom[120][7] = 16'hFFF3;
        rom[120][8] = 16'h0008;
        rom[120][9] = 16'hFFFE;
        rom[120][10] = 16'h0002;
        rom[120][11] = 16'h0016;
        rom[120][12] = 16'h0007;
        rom[120][13] = 16'h0007;
        rom[120][14] = 16'hFFFB;
        rom[120][15] = 16'h001B;
        rom[120][16] = 16'h0000;
        rom[120][17] = 16'h001B;
        rom[120][18] = 16'hFFDC;
        rom[120][19] = 16'h000F;
        rom[120][20] = 16'hFFE2;
        rom[120][21] = 16'h0017;
        rom[120][22] = 16'h0013;
        rom[120][23] = 16'hFFEB;
        rom[120][24] = 16'h0015;
        rom[120][25] = 16'hFFFE;
        rom[120][26] = 16'hFFD7;
        rom[120][27] = 16'hFFE9;
        rom[120][28] = 16'hFFF0;
        rom[120][29] = 16'h0001;
        rom[120][30] = 16'hFFF2;
        rom[120][31] = 16'h002C;
        rom[120][32] = 16'hFFF0;
        rom[120][33] = 16'h0011;
        rom[120][34] = 16'h0024;
        rom[120][35] = 16'h0020;
        rom[120][36] = 16'h001E;
        rom[120][37] = 16'h000B;
        rom[120][38] = 16'h0025;
        rom[120][39] = 16'h0001;
        rom[120][40] = 16'hFFFD;
        rom[120][41] = 16'h0015;
        rom[120][42] = 16'hFFD2;
        rom[120][43] = 16'hFFC5;
        rom[120][44] = 16'h0019;
        rom[120][45] = 16'h0011;
        rom[120][46] = 16'hFFE4;
        rom[120][47] = 16'hFFE3;
        rom[120][48] = 16'hFFFB;
        rom[120][49] = 16'h0017;
        rom[120][50] = 16'hFFF4;
        rom[120][51] = 16'h0011;
        rom[120][52] = 16'hFFC8;
        rom[120][53] = 16'hFFD0;
        rom[120][54] = 16'h000D;
        rom[120][55] = 16'hFFD7;
        rom[120][56] = 16'h001E;
        rom[120][57] = 16'hFFD1;
        rom[120][58] = 16'h0008;
        rom[120][59] = 16'hFFF6;
        rom[120][60] = 16'h0002;
        rom[120][61] = 16'h000B;
        rom[120][62] = 16'hFFE8;
        rom[120][63] = 16'hFFF7;
        rom[120][64] = 16'hFFF1;
        rom[120][65] = 16'h0009;
        rom[120][66] = 16'hFFED;
        rom[120][67] = 16'hFFBF;
        rom[120][68] = 16'h0029;
        rom[120][69] = 16'hFFEF;
        rom[120][70] = 16'h0024;
        rom[120][71] = 16'hFFD0;
        rom[120][72] = 16'h0003;
        rom[120][73] = 16'h001C;
        rom[120][74] = 16'hFFFB;
        rom[120][75] = 16'h001C;
        rom[120][76] = 16'h000E;
        rom[120][77] = 16'hFFEF;
        rom[120][78] = 16'h0006;
        rom[120][79] = 16'hFFD6;
        rom[120][80] = 16'hFFC8;
        rom[120][81] = 16'h0011;
        rom[120][82] = 16'hFFD7;
        rom[120][83] = 16'h002B;
        rom[120][84] = 16'h0000;
        rom[120][85] = 16'hFFF4;
        rom[120][86] = 16'h0003;
        rom[120][87] = 16'hFFDA;
        rom[120][88] = 16'h001B;
        rom[120][89] = 16'h000C;
        rom[120][90] = 16'hFFBF;
        rom[120][91] = 16'hFFE3;
        rom[120][92] = 16'h0011;
        rom[120][93] = 16'h000E;
        rom[120][94] = 16'hFFF1;
        rom[120][95] = 16'hFFD9;
        rom[120][96] = 16'h0005;
        rom[120][97] = 16'hFFD2;
        rom[120][98] = 16'h0014;
        rom[120][99] = 16'h0009;
        rom[120][100] = 16'hFFB8;
        rom[120][101] = 16'hFFA2;
        rom[120][102] = 16'hFFEB;
        rom[120][103] = 16'hFFF3;
        rom[120][104] = 16'hFFE4;
        rom[120][105] = 16'h000D;
        rom[120][106] = 16'hFFE1;
        rom[120][107] = 16'h000A;
        rom[120][108] = 16'hFFE2;
        rom[120][109] = 16'h000B;
        rom[120][110] = 16'hFFEA;
        rom[120][111] = 16'h0024;
        rom[120][112] = 16'hFFF5;
        rom[120][113] = 16'hFFEC;
        rom[120][114] = 16'h0014;
        rom[120][115] = 16'h002D;
        rom[120][116] = 16'h000C;
        rom[120][117] = 16'h000F;
        rom[120][118] = 16'hFFAF;
        rom[120][119] = 16'h0022;
        rom[120][120] = 16'h0007;
        rom[120][121] = 16'h0008;
        rom[120][122] = 16'hFFFD;
        rom[120][123] = 16'h000A;
        rom[120][124] = 16'h0000;
        rom[120][125] = 16'hFFD1;
        rom[120][126] = 16'hFFDF;
        rom[120][127] = 16'hFFD9;
        rom[121][0] = 16'h0004;
        rom[121][1] = 16'hFFF7;
        rom[121][2] = 16'hFFE9;
        rom[121][3] = 16'h000B;
        rom[121][4] = 16'hFFD5;
        rom[121][5] = 16'hFFED;
        rom[121][6] = 16'hFFFA;
        rom[121][7] = 16'hFFFD;
        rom[121][8] = 16'hFFC9;
        rom[121][9] = 16'h0007;
        rom[121][10] = 16'hFFE0;
        rom[121][11] = 16'hFFD7;
        rom[121][12] = 16'hFFDC;
        rom[121][13] = 16'h000E;
        rom[121][14] = 16'h0006;
        rom[121][15] = 16'hFFF4;
        rom[121][16] = 16'hFFF2;
        rom[121][17] = 16'hFFD0;
        rom[121][18] = 16'h0029;
        rom[121][19] = 16'hFFEE;
        rom[121][20] = 16'hFFFC;
        rom[121][21] = 16'h0018;
        rom[121][22] = 16'hFFC8;
        rom[121][23] = 16'hFFE1;
        rom[121][24] = 16'h001B;
        rom[121][25] = 16'h0011;
        rom[121][26] = 16'hFFEF;
        rom[121][27] = 16'hFFDA;
        rom[121][28] = 16'hFFEF;
        rom[121][29] = 16'h0000;
        rom[121][30] = 16'h002A;
        rom[121][31] = 16'h0002;
        rom[121][32] = 16'hFFD0;
        rom[121][33] = 16'h0012;
        rom[121][34] = 16'hFFCA;
        rom[121][35] = 16'h0016;
        rom[121][36] = 16'h000A;
        rom[121][37] = 16'h0007;
        rom[121][38] = 16'hFFE5;
        rom[121][39] = 16'h0031;
        rom[121][40] = 16'h001C;
        rom[121][41] = 16'hFFEF;
        rom[121][42] = 16'hFFE6;
        rom[121][43] = 16'hFFFE;
        rom[121][44] = 16'h002A;
        rom[121][45] = 16'hFFEB;
        rom[121][46] = 16'hFFEA;
        rom[121][47] = 16'hFFCA;
        rom[121][48] = 16'h0006;
        rom[121][49] = 16'hFFF1;
        rom[121][50] = 16'hFFFA;
        rom[121][51] = 16'h0028;
        rom[121][52] = 16'h0013;
        rom[121][53] = 16'h0020;
        rom[121][54] = 16'hFFC0;
        rom[121][55] = 16'h0007;
        rom[121][56] = 16'h000A;
        rom[121][57] = 16'hFFE2;
        rom[121][58] = 16'hFFC9;
        rom[121][59] = 16'hFFB5;
        rom[121][60] = 16'h000D;
        rom[121][61] = 16'h000C;
        rom[121][62] = 16'hFFEA;
        rom[121][63] = 16'hFFF4;
        rom[121][64] = 16'h0016;
        rom[121][65] = 16'h000A;
        rom[121][66] = 16'h000F;
        rom[121][67] = 16'hFFE6;
        rom[121][68] = 16'h0015;
        rom[121][69] = 16'h0004;
        rom[121][70] = 16'hFFF9;
        rom[121][71] = 16'h0013;
        rom[121][72] = 16'hFFE7;
        rom[121][73] = 16'h0000;
        rom[121][74] = 16'hFFF9;
        rom[121][75] = 16'h0025;
        rom[121][76] = 16'h001E;
        rom[121][77] = 16'h0066;
        rom[121][78] = 16'h0004;
        rom[121][79] = 16'h001F;
        rom[121][80] = 16'hFFD2;
        rom[121][81] = 16'hFFD9;
        rom[121][82] = 16'hFFE4;
        rom[121][83] = 16'h001D;
        rom[121][84] = 16'hFFF2;
        rom[121][85] = 16'hFFDC;
        rom[121][86] = 16'h0026;
        rom[121][87] = 16'hFFBA;
        rom[121][88] = 16'h0006;
        rom[121][89] = 16'hFFB0;
        rom[121][90] = 16'hFFFC;
        rom[121][91] = 16'hFFFA;
        rom[121][92] = 16'h0014;
        rom[121][93] = 16'hFFFD;
        rom[121][94] = 16'hFFD5;
        rom[121][95] = 16'h0007;
        rom[121][96] = 16'hFFCC;
        rom[121][97] = 16'hFFDC;
        rom[121][98] = 16'h0029;
        rom[121][99] = 16'hFFF5;
        rom[121][100] = 16'hFFE5;
        rom[121][101] = 16'h002E;
        rom[121][102] = 16'h0006;
        rom[121][103] = 16'hFFF3;
        rom[121][104] = 16'h0027;
        rom[121][105] = 16'h0014;
        rom[121][106] = 16'h0006;
        rom[121][107] = 16'hFFC3;
        rom[121][108] = 16'hFFED;
        rom[121][109] = 16'h0017;
        rom[121][110] = 16'hFFCA;
        rom[121][111] = 16'hFFF9;
        rom[121][112] = 16'hFFF9;
        rom[121][113] = 16'h001F;
        rom[121][114] = 16'h0002;
        rom[121][115] = 16'h0004;
        rom[121][116] = 16'hFFFE;
        rom[121][117] = 16'h0005;
        rom[121][118] = 16'hFFD6;
        rom[121][119] = 16'hFFE0;
        rom[121][120] = 16'h0022;
        rom[121][121] = 16'hFFDC;
        rom[121][122] = 16'hFFCC;
        rom[121][123] = 16'h0013;
        rom[121][124] = 16'hFFCD;
        rom[121][125] = 16'hFFF1;
        rom[121][126] = 16'hFFC9;
        rom[121][127] = 16'hFFF0;
        rom[122][0] = 16'h000A;
        rom[122][1] = 16'h0008;
        rom[122][2] = 16'hFFC3;
        rom[122][3] = 16'hFFC8;
        rom[122][4] = 16'hFFF5;
        rom[122][5] = 16'hFFF4;
        rom[122][6] = 16'h000B;
        rom[122][7] = 16'h000D;
        rom[122][8] = 16'h0005;
        rom[122][9] = 16'hFFCC;
        rom[122][10] = 16'hFFFD;
        rom[122][11] = 16'hFFD4;
        rom[122][12] = 16'hFFF4;
        rom[122][13] = 16'hFFDF;
        rom[122][14] = 16'hFFF9;
        rom[122][15] = 16'h0009;
        rom[122][16] = 16'h0008;
        rom[122][17] = 16'hFFB8;
        rom[122][18] = 16'hFFD2;
        rom[122][19] = 16'h0011;
        rom[122][20] = 16'h0011;
        rom[122][21] = 16'hFFDC;
        rom[122][22] = 16'hFFC8;
        rom[122][23] = 16'hFFC4;
        rom[122][24] = 16'hFFEE;
        rom[122][25] = 16'h001D;
        rom[122][26] = 16'hFFF7;
        rom[122][27] = 16'h0007;
        rom[122][28] = 16'h001E;
        rom[122][29] = 16'h0019;
        rom[122][30] = 16'h0001;
        rom[122][31] = 16'h001B;
        rom[122][32] = 16'hFFD2;
        rom[122][33] = 16'hFFBA;
        rom[122][34] = 16'hFFF6;
        rom[122][35] = 16'h000C;
        rom[122][36] = 16'h001B;
        rom[122][37] = 16'hFFF4;
        rom[122][38] = 16'hFFDC;
        rom[122][39] = 16'h0013;
        rom[122][40] = 16'h0000;
        rom[122][41] = 16'h0005;
        rom[122][42] = 16'hFFEF;
        rom[122][43] = 16'hFFCE;
        rom[122][44] = 16'h0010;
        rom[122][45] = 16'hFFF4;
        rom[122][46] = 16'h0015;
        rom[122][47] = 16'hFFF1;
        rom[122][48] = 16'h0013;
        rom[122][49] = 16'h000C;
        rom[122][50] = 16'hFFC3;
        rom[122][51] = 16'hFFD4;
        rom[122][52] = 16'hFFA2;
        rom[122][53] = 16'hFFAE;
        rom[122][54] = 16'h0001;
        rom[122][55] = 16'hFFF4;
        rom[122][56] = 16'hFFF8;
        rom[122][57] = 16'hFFF9;
        rom[122][58] = 16'h0002;
        rom[122][59] = 16'h000D;
        rom[122][60] = 16'h0007;
        rom[122][61] = 16'h001E;
        rom[122][62] = 16'h0003;
        rom[122][63] = 16'h0013;
        rom[122][64] = 16'h0015;
        rom[122][65] = 16'h0000;
        rom[122][66] = 16'hFFED;
        rom[122][67] = 16'hFFD6;
        rom[122][68] = 16'hFFE9;
        rom[122][69] = 16'hFFFD;
        rom[122][70] = 16'hFFA1;
        rom[122][71] = 16'hFFC1;
        rom[122][72] = 16'h0011;
        rom[122][73] = 16'hFFFF;
        rom[122][74] = 16'h001C;
        rom[122][75] = 16'hFFD0;
        rom[122][76] = 16'hFFEC;
        rom[122][77] = 16'hFFCB;
        rom[122][78] = 16'h0002;
        rom[122][79] = 16'h0018;
        rom[122][80] = 16'h0009;
        rom[122][81] = 16'hFFFB;
        rom[122][82] = 16'h0012;
        rom[122][83] = 16'h001B;
        rom[122][84] = 16'h0013;
        rom[122][85] = 16'hFFFC;
        rom[122][86] = 16'h002E;
        rom[122][87] = 16'hFFCC;
        rom[122][88] = 16'h0011;
        rom[122][89] = 16'hFFFA;
        rom[122][90] = 16'h000C;
        rom[122][91] = 16'hFFFB;
        rom[122][92] = 16'hFFD1;
        rom[122][93] = 16'h000A;
        rom[122][94] = 16'hFFBA;
        rom[122][95] = 16'h0012;
        rom[122][96] = 16'h0002;
        rom[122][97] = 16'h0008;
        rom[122][98] = 16'h0010;
        rom[122][99] = 16'h0002;
        rom[122][100] = 16'h0013;
        rom[122][101] = 16'h001A;
        rom[122][102] = 16'hFFF6;
        rom[122][103] = 16'hFFCF;
        rom[122][104] = 16'hFFED;
        rom[122][105] = 16'hFFE1;
        rom[122][106] = 16'h0007;
        rom[122][107] = 16'hFFE0;
        rom[122][108] = 16'h000C;
        rom[122][109] = 16'h000B;
        rom[122][110] = 16'h0017;
        rom[122][111] = 16'h0021;
        rom[122][112] = 16'h0001;
        rom[122][113] = 16'hFFF4;
        rom[122][114] = 16'hFFF9;
        rom[122][115] = 16'h001D;
        rom[122][116] = 16'hFFFF;
        rom[122][117] = 16'h001F;
        rom[122][118] = 16'hFFE5;
        rom[122][119] = 16'hFFD1;
        rom[122][120] = 16'hFFFE;
        rom[122][121] = 16'hFFF1;
        rom[122][122] = 16'hFFC3;
        rom[122][123] = 16'hFFAE;
        rom[122][124] = 16'hFFEC;
        rom[122][125] = 16'hFFC5;
        rom[122][126] = 16'hFFC8;
        rom[122][127] = 16'hFFEF;
        rom[123][0] = 16'h0018;
        rom[123][1] = 16'h0002;
        rom[123][2] = 16'h0004;
        rom[123][3] = 16'hFFEA;
        rom[123][4] = 16'hFFFF;
        rom[123][5] = 16'hFFF4;
        rom[123][6] = 16'hFFF1;
        rom[123][7] = 16'h001A;
        rom[123][8] = 16'h0006;
        rom[123][9] = 16'hFFEB;
        rom[123][10] = 16'hFFA9;
        rom[123][11] = 16'h0000;
        rom[123][12] = 16'hFFF2;
        rom[123][13] = 16'hFFD0;
        rom[123][14] = 16'hFFDD;
        rom[123][15] = 16'h0007;
        rom[123][16] = 16'hFFD2;
        rom[123][17] = 16'hFFC9;
        rom[123][18] = 16'h0011;
        rom[123][19] = 16'hFFC4;
        rom[123][20] = 16'hFFE5;
        rom[123][21] = 16'h0048;
        rom[123][22] = 16'hFFEB;
        rom[123][23] = 16'hFFEA;
        rom[123][24] = 16'h0019;
        rom[123][25] = 16'hFFCD;
        rom[123][26] = 16'h0007;
        rom[123][27] = 16'hFFFE;
        rom[123][28] = 16'h000C;
        rom[123][29] = 16'hFFC4;
        rom[123][30] = 16'h0014;
        rom[123][31] = 16'hFFFA;
        rom[123][32] = 16'hFFD8;
        rom[123][33] = 16'h0022;
        rom[123][34] = 16'hFFE0;
        rom[123][35] = 16'hFFEF;
        rom[123][36] = 16'hFFEF;
        rom[123][37] = 16'hFFF7;
        rom[123][38] = 16'h0005;
        rom[123][39] = 16'h002E;
        rom[123][40] = 16'hFFB2;
        rom[123][41] = 16'hFFCB;
        rom[123][42] = 16'h0001;
        rom[123][43] = 16'hFFD2;
        rom[123][44] = 16'hFFD7;
        rom[123][45] = 16'h0011;
        rom[123][46] = 16'h0000;
        rom[123][47] = 16'h0007;
        rom[123][48] = 16'hFFC6;
        rom[123][49] = 16'hFFEC;
        rom[123][50] = 16'h0008;
        rom[123][51] = 16'h0015;
        rom[123][52] = 16'hFFF8;
        rom[123][53] = 16'hFFDF;
        rom[123][54] = 16'h001B;
        rom[123][55] = 16'h001D;
        rom[123][56] = 16'hFFE1;
        rom[123][57] = 16'hFFC8;
        rom[123][58] = 16'h0007;
        rom[123][59] = 16'hFFDA;
        rom[123][60] = 16'h0033;
        rom[123][61] = 16'hFFB8;
        rom[123][62] = 16'hFFFA;
        rom[123][63] = 16'h0011;
        rom[123][64] = 16'hFFF4;
        rom[123][65] = 16'h001A;
        rom[123][66] = 16'h0005;
        rom[123][67] = 16'hFFE6;
        rom[123][68] = 16'h0014;
        rom[123][69] = 16'h000C;
        rom[123][70] = 16'h0016;
        rom[123][71] = 16'h000F;
        rom[123][72] = 16'h0014;
        rom[123][73] = 16'h0011;
        rom[123][74] = 16'h000D;
        rom[123][75] = 16'h0038;
        rom[123][76] = 16'hFFEA;
        rom[123][77] = 16'h0005;
        rom[123][78] = 16'h0026;
        rom[123][79] = 16'hFFF8;
        rom[123][80] = 16'hFFFA;
        rom[123][81] = 16'h001B;
        rom[123][82] = 16'hFFEB;
        rom[123][83] = 16'h000D;
        rom[123][84] = 16'hFFFD;
        rom[123][85] = 16'h0004;
        rom[123][86] = 16'hFFEC;
        rom[123][87] = 16'hFFEA;
        rom[123][88] = 16'hFFEA;
        rom[123][89] = 16'h0012;
        rom[123][90] = 16'hFFD8;
        rom[123][91] = 16'hFFD7;
        rom[123][92] = 16'h004D;
        rom[123][93] = 16'h001B;
        rom[123][94] = 16'hFFF0;
        rom[123][95] = 16'h002C;
        rom[123][96] = 16'hFFBF;
        rom[123][97] = 16'hFFAC;
        rom[123][98] = 16'hFFE0;
        rom[123][99] = 16'h0009;
        rom[123][100] = 16'h0034;
        rom[123][101] = 16'h002C;
        rom[123][102] = 16'h0000;
        rom[123][103] = 16'hFFEE;
        rom[123][104] = 16'h0011;
        rom[123][105] = 16'hFFBA;
        rom[123][106] = 16'h000E;
        rom[123][107] = 16'hFFFE;
        rom[123][108] = 16'hFFD7;
        rom[123][109] = 16'h0016;
        rom[123][110] = 16'hFFF9;
        rom[123][111] = 16'h000E;
        rom[123][112] = 16'hFFFF;
        rom[123][113] = 16'h0004;
        rom[123][114] = 16'hFFEA;
        rom[123][115] = 16'hFFF0;
        rom[123][116] = 16'h0005;
        rom[123][117] = 16'hFFD4;
        rom[123][118] = 16'h0017;
        rom[123][119] = 16'h0020;
        rom[123][120] = 16'h000C;
        rom[123][121] = 16'hFFFE;
        rom[123][122] = 16'hFFF3;
        rom[123][123] = 16'h0012;
        rom[123][124] = 16'hFFF3;
        rom[123][125] = 16'h0023;
        rom[123][126] = 16'hFFB5;
        rom[123][127] = 16'hFFBB;
        rom[124][0] = 16'hFFE6;
        rom[124][1] = 16'h0011;
        rom[124][2] = 16'h001A;
        rom[124][3] = 16'h001C;
        rom[124][4] = 16'hFFBB;
        rom[124][5] = 16'h0018;
        rom[124][6] = 16'h0007;
        rom[124][7] = 16'hFFF1;
        rom[124][8] = 16'h000D;
        rom[124][9] = 16'hFFF2;
        rom[124][10] = 16'hFFC1;
        rom[124][11] = 16'h0027;
        rom[124][12] = 16'hFFA3;
        rom[124][13] = 16'hFFF9;
        rom[124][14] = 16'h0002;
        rom[124][15] = 16'hFFE9;
        rom[124][16] = 16'hFFE1;
        rom[124][17] = 16'h001C;
        rom[124][18] = 16'h000A;
        rom[124][19] = 16'hFFE9;
        rom[124][20] = 16'hFFEA;
        rom[124][21] = 16'h0007;
        rom[124][22] = 16'hFFFF;
        rom[124][23] = 16'h0003;
        rom[124][24] = 16'hFFB1;
        rom[124][25] = 16'hFFFA;
        rom[124][26] = 16'h0008;
        rom[124][27] = 16'hFFB3;
        rom[124][28] = 16'hFFE9;
        rom[124][29] = 16'h0009;
        rom[124][30] = 16'hFFCF;
        rom[124][31] = 16'h0019;
        rom[124][32] = 16'h003F;
        rom[124][33] = 16'hFFC3;
        rom[124][34] = 16'hFFCA;
        rom[124][35] = 16'h0009;
        rom[124][36] = 16'h0010;
        rom[124][37] = 16'h001D;
        rom[124][38] = 16'hFFF9;
        rom[124][39] = 16'hFFF1;
        rom[124][40] = 16'h000C;
        rom[124][41] = 16'hFFE5;
        rom[124][42] = 16'hFFEB;
        rom[124][43] = 16'hFFE0;
        rom[124][44] = 16'hFFDB;
        rom[124][45] = 16'h0018;
        rom[124][46] = 16'h0006;
        rom[124][47] = 16'h0005;
        rom[124][48] = 16'hFFEF;
        rom[124][49] = 16'hFFD4;
        rom[124][50] = 16'hFFF4;
        rom[124][51] = 16'h0002;
        rom[124][52] = 16'h0005;
        rom[124][53] = 16'h0004;
        rom[124][54] = 16'h0015;
        rom[124][55] = 16'hFFDC;
        rom[124][56] = 16'h0009;
        rom[124][57] = 16'hFFE9;
        rom[124][58] = 16'h0002;
        rom[124][59] = 16'h0028;
        rom[124][60] = 16'hFFD8;
        rom[124][61] = 16'hFFD2;
        rom[124][62] = 16'hFFFA;
        rom[124][63] = 16'h001A;
        rom[124][64] = 16'hFFEE;
        rom[124][65] = 16'hFFF1;
        rom[124][66] = 16'h0002;
        rom[124][67] = 16'h000C;
        rom[124][68] = 16'h002F;
        rom[124][69] = 16'hFFD2;
        rom[124][70] = 16'hFFE3;
        rom[124][71] = 16'h0030;
        rom[124][72] = 16'hFFE2;
        rom[124][73] = 16'h0014;
        rom[124][74] = 16'h000B;
        rom[124][75] = 16'hFFAA;
        rom[124][76] = 16'hFFEB;
        rom[124][77] = 16'hFFE3;
        rom[124][78] = 16'h0024;
        rom[124][79] = 16'hFFF1;
        rom[124][80] = 16'h0020;
        rom[124][81] = 16'h0029;
        rom[124][82] = 16'h0013;
        rom[124][83] = 16'hFFDD;
        rom[124][84] = 16'h0000;
        rom[124][85] = 16'hFFE6;
        rom[124][86] = 16'h000E;
        rom[124][87] = 16'h000E;
        rom[124][88] = 16'hFFF8;
        rom[124][89] = 16'h0005;
        rom[124][90] = 16'h001F;
        rom[124][91] = 16'hFFF5;
        rom[124][92] = 16'hFFB9;
        rom[124][93] = 16'h0008;
        rom[124][94] = 16'h0010;
        rom[124][95] = 16'h001C;
        rom[124][96] = 16'hFFEC;
        rom[124][97] = 16'hFFD9;
        rom[124][98] = 16'hFFC2;
        rom[124][99] = 16'h0001;
        rom[124][100] = 16'hFFD6;
        rom[124][101] = 16'hFFEA;
        rom[124][102] = 16'hFFBA;
        rom[124][103] = 16'hFFCA;
        rom[124][104] = 16'h0026;
        rom[124][105] = 16'hFFF8;
        rom[124][106] = 16'h0011;
        rom[124][107] = 16'h002D;
        rom[124][108] = 16'hFFD2;
        rom[124][109] = 16'h0009;
        rom[124][110] = 16'hFFE9;
        rom[124][111] = 16'hFFF9;
        rom[124][112] = 16'hFFE5;
        rom[124][113] = 16'hFFB8;
        rom[124][114] = 16'hFFBF;
        rom[124][115] = 16'h0000;
        rom[124][116] = 16'hFFD1;
        rom[124][117] = 16'hFFCD;
        rom[124][118] = 16'hFFED;
        rom[124][119] = 16'h0000;
        rom[124][120] = 16'h0005;
        rom[124][121] = 16'hFFF4;
        rom[124][122] = 16'h0015;
        rom[124][123] = 16'hFFD2;
        rom[124][124] = 16'h0009;
        rom[124][125] = 16'h0009;
        rom[124][126] = 16'hFFF7;
        rom[124][127] = 16'h0007;
        rom[125][0] = 16'hFFF5;
        rom[125][1] = 16'h0020;
        rom[125][2] = 16'h0006;
        rom[125][3] = 16'h0002;
        rom[125][4] = 16'hFFDF;
        rom[125][5] = 16'h0031;
        rom[125][6] = 16'hFFDE;
        rom[125][7] = 16'h0002;
        rom[125][8] = 16'h0001;
        rom[125][9] = 16'h0027;
        rom[125][10] = 16'hFFD8;
        rom[125][11] = 16'hFFB5;
        rom[125][12] = 16'hFFE6;
        rom[125][13] = 16'hFFCA;
        rom[125][14] = 16'h001A;
        rom[125][15] = 16'h0003;
        rom[125][16] = 16'hFFD2;
        rom[125][17] = 16'hFFD3;
        rom[125][18] = 16'hFFE5;
        rom[125][19] = 16'hFFFC;
        rom[125][20] = 16'hFFEF;
        rom[125][21] = 16'hFFF4;
        rom[125][22] = 16'hFFFC;
        rom[125][23] = 16'h0012;
        rom[125][24] = 16'h0014;
        rom[125][25] = 16'hFFEA;
        rom[125][26] = 16'hFFE1;
        rom[125][27] = 16'hFFBB;
        rom[125][28] = 16'hFFC2;
        rom[125][29] = 16'hFFEF;
        rom[125][30] = 16'hFFEE;
        rom[125][31] = 16'hFFF2;
        rom[125][32] = 16'hFFEA;
        rom[125][33] = 16'h000B;
        rom[125][34] = 16'hFFEA;
        rom[125][35] = 16'hFFD5;
        rom[125][36] = 16'hFFFB;
        rom[125][37] = 16'hFFE3;
        rom[125][38] = 16'hFFFC;
        rom[125][39] = 16'h0033;
        rom[125][40] = 16'hFFDD;
        rom[125][41] = 16'h0005;
        rom[125][42] = 16'h000C;
        rom[125][43] = 16'hFFEF;
        rom[125][44] = 16'hFFE4;
        rom[125][45] = 16'hFFF6;
        rom[125][46] = 16'h000A;
        rom[125][47] = 16'h0009;
        rom[125][48] = 16'h0005;
        rom[125][49] = 16'hFFFE;
        rom[125][50] = 16'h0035;
        rom[125][51] = 16'hFFEA;
        rom[125][52] = 16'h0013;
        rom[125][53] = 16'h001F;
        rom[125][54] = 16'hFFF2;
        rom[125][55] = 16'h0017;
        rom[125][56] = 16'hFFD1;
        rom[125][57] = 16'h0005;
        rom[125][58] = 16'h0020;
        rom[125][59] = 16'hFFC9;
        rom[125][60] = 16'h0005;
        rom[125][61] = 16'hFFE2;
        rom[125][62] = 16'h0002;
        rom[125][63] = 16'h000D;
        rom[125][64] = 16'hFFCD;
        rom[125][65] = 16'h000C;
        rom[125][66] = 16'h0011;
        rom[125][67] = 16'hFFFF;
        rom[125][68] = 16'hFFDC;
        rom[125][69] = 16'h0007;
        rom[125][70] = 16'h0028;
        rom[125][71] = 16'h0002;
        rom[125][72] = 16'hFFCB;
        rom[125][73] = 16'hFFED;
        rom[125][74] = 16'hFFE3;
        rom[125][75] = 16'hFFF6;
        rom[125][76] = 16'hFFFC;
        rom[125][77] = 16'hFFF9;
        rom[125][78] = 16'h000F;
        rom[125][79] = 16'hFFF9;
        rom[125][80] = 16'h000A;
        rom[125][81] = 16'h0002;
        rom[125][82] = 16'h001A;
        rom[125][83] = 16'h0010;
        rom[125][84] = 16'hFFFA;
        rom[125][85] = 16'h0020;
        rom[125][86] = 16'hFFE2;
        rom[125][87] = 16'h0007;
        rom[125][88] = 16'hFFDF;
        rom[125][89] = 16'hFFFE;
        rom[125][90] = 16'hFFD8;
        rom[125][91] = 16'h001B;
        rom[125][92] = 16'h0009;
        rom[125][93] = 16'hFFED;
        rom[125][94] = 16'h000E;
        rom[125][95] = 16'h0026;
        rom[125][96] = 16'hFFFB;
        rom[125][97] = 16'h000F;
        rom[125][98] = 16'hFFB6;
        rom[125][99] = 16'h0012;
        rom[125][100] = 16'hFFD4;
        rom[125][101] = 16'hFFD2;
        rom[125][102] = 16'hFFF5;
        rom[125][103] = 16'hFFD6;
        rom[125][104] = 16'hFFD9;
        rom[125][105] = 16'h001B;
        rom[125][106] = 16'hFFFF;
        rom[125][107] = 16'hFFF9;
        rom[125][108] = 16'hFFF3;
        rom[125][109] = 16'hFFDB;
        rom[125][110] = 16'hFFD7;
        rom[125][111] = 16'hFFFE;
        rom[125][112] = 16'hFFFA;
        rom[125][113] = 16'h002E;
        rom[125][114] = 16'hFFDC;
        rom[125][115] = 16'h000B;
        rom[125][116] = 16'h0011;
        rom[125][117] = 16'h002C;
        rom[125][118] = 16'h000A;
        rom[125][119] = 16'h0001;
        rom[125][120] = 16'hFFEF;
        rom[125][121] = 16'h0030;
        rom[125][122] = 16'hFFFD;
        rom[125][123] = 16'h0017;
        rom[125][124] = 16'hFFF2;
        rom[125][125] = 16'hFFF0;
        rom[125][126] = 16'h0005;
        rom[125][127] = 16'hFFCC;
        rom[126][0] = 16'h0018;
        rom[126][1] = 16'h0017;
        rom[126][2] = 16'h0014;
        rom[126][3] = 16'h0007;
        rom[126][4] = 16'hFFD6;
        rom[126][5] = 16'h0003;
        rom[126][6] = 16'hFFF9;
        rom[126][7] = 16'h0011;
        rom[126][8] = 16'h0021;
        rom[126][9] = 16'h0021;
        rom[126][10] = 16'hFFDE;
        rom[126][11] = 16'hFFFA;
        rom[126][12] = 16'h0033;
        rom[126][13] = 16'h0012;
        rom[126][14] = 16'hFFF4;
        rom[126][15] = 16'h0001;
        rom[126][16] = 16'hFFD7;
        rom[126][17] = 16'h0020;
        rom[126][18] = 16'h0005;
        rom[126][19] = 16'h0010;
        rom[126][20] = 16'hFFFE;
        rom[126][21] = 16'h0007;
        rom[126][22] = 16'h001C;
        rom[126][23] = 16'h0004;
        rom[126][24] = 16'h0018;
        rom[126][25] = 16'h0024;
        rom[126][26] = 16'hFFF8;
        rom[126][27] = 16'h0007;
        rom[126][28] = 16'hFFAB;
        rom[126][29] = 16'hFFF4;
        rom[126][30] = 16'hFFDC;
        rom[126][31] = 16'hFFFE;
        rom[126][32] = 16'h0007;
        rom[126][33] = 16'h0007;
        rom[126][34] = 16'h0007;
        rom[126][35] = 16'h0007;
        rom[126][36] = 16'h001F;
        rom[126][37] = 16'h0009;
        rom[126][38] = 16'h0036;
        rom[126][39] = 16'h0029;
        rom[126][40] = 16'hFFFC;
        rom[126][41] = 16'h0007;
        rom[126][42] = 16'h0021;
        rom[126][43] = 16'hFFC5;
        rom[126][44] = 16'hFFF4;
        rom[126][45] = 16'hFFFC;
        rom[126][46] = 16'h0020;
        rom[126][47] = 16'h002B;
        rom[126][48] = 16'h0012;
        rom[126][49] = 16'h0003;
        rom[126][50] = 16'h0019;
        rom[126][51] = 16'h0001;
        rom[126][52] = 16'h005C;
        rom[126][53] = 16'hFFFB;
        rom[126][54] = 16'hFFE2;
        rom[126][55] = 16'hFFFA;
        rom[126][56] = 16'hFFFE;
        rom[126][57] = 16'h0009;
        rom[126][58] = 16'h0017;
        rom[126][59] = 16'hFFFA;
        rom[126][60] = 16'hFFA6;
        rom[126][61] = 16'hFFF4;
        rom[126][62] = 16'h0003;
        rom[126][63] = 16'h000F;
        rom[126][64] = 16'hFFF8;
        rom[126][65] = 16'hFFF5;
        rom[126][66] = 16'h0013;
        rom[126][67] = 16'h0007;
        rom[126][68] = 16'hFFDD;
        rom[126][69] = 16'hFFEF;
        rom[126][70] = 16'h0023;
        rom[126][71] = 16'hFFA8;
        rom[126][72] = 16'h002F;
        rom[126][73] = 16'hFFF0;
        rom[126][74] = 16'hFFF7;
        rom[126][75] = 16'h0006;
        rom[126][76] = 16'h000A;
        rom[126][77] = 16'hFFBD;
        rom[126][78] = 16'hFFD2;
        rom[126][79] = 16'hFFEE;
        rom[126][80] = 16'h0001;
        rom[126][81] = 16'hFFD6;
        rom[126][82] = 16'hFFFB;
        rom[126][83] = 16'h001E;
        rom[126][84] = 16'h0007;
        rom[126][85] = 16'h0019;
        rom[126][86] = 16'h000E;
        rom[126][87] = 16'hFFCC;
        rom[126][88] = 16'hFFEF;
        rom[126][89] = 16'hFFE9;
        rom[126][90] = 16'hFFEA;
        rom[126][91] = 16'hFFD1;
        rom[126][92] = 16'h0008;
        rom[126][93] = 16'hFFC5;
        rom[126][94] = 16'hFFF0;
        rom[126][95] = 16'h001C;
        rom[126][96] = 16'hFFDD;
        rom[126][97] = 16'hFFD3;
        rom[126][98] = 16'hFFB5;
        rom[126][99] = 16'hFFD8;
        rom[126][100] = 16'hFFA9;
        rom[126][101] = 16'hFFFA;
        rom[126][102] = 16'h0004;
        rom[126][103] = 16'h0017;
        rom[126][104] = 16'hFFEB;
        rom[126][105] = 16'h0010;
        rom[126][106] = 16'h0008;
        rom[126][107] = 16'hFFF4;
        rom[126][108] = 16'hFFA2;
        rom[126][109] = 16'h000F;
        rom[126][110] = 16'h002F;
        rom[126][111] = 16'hFFDD;
        rom[126][112] = 16'h0029;
        rom[126][113] = 16'h0025;
        rom[126][114] = 16'hFFE9;
        rom[126][115] = 16'hFFFD;
        rom[126][116] = 16'h0011;
        rom[126][117] = 16'h0020;
        rom[126][118] = 16'h0019;
        rom[126][119] = 16'h0029;
        rom[126][120] = 16'h0016;
        rom[126][121] = 16'h001A;
        rom[126][122] = 16'hFFD7;
        rom[126][123] = 16'h0024;
        rom[126][124] = 16'hFFE8;
        rom[126][125] = 16'hFFD3;
        rom[126][126] = 16'hFFEF;
        rom[126][127] = 16'hFFF3;
        rom[127][0] = 16'h0028;
        rom[127][1] = 16'hFFF0;
        rom[127][2] = 16'hFFDB;
        rom[127][3] = 16'h0011;
        rom[127][4] = 16'hFFD7;
        rom[127][5] = 16'hFFE4;
        rom[127][6] = 16'hFFAA;
        rom[127][7] = 16'h001F;
        rom[127][8] = 16'hFFD5;
        rom[127][9] = 16'hFFA2;
        rom[127][10] = 16'hFFCF;
        rom[127][11] = 16'hFFF9;
        rom[127][12] = 16'h0007;
        rom[127][13] = 16'hFFFE;
        rom[127][14] = 16'hFFFB;
        rom[127][15] = 16'h000C;
        rom[127][16] = 16'hFFCB;
        rom[127][17] = 16'h0011;
        rom[127][18] = 16'hFFDF;
        rom[127][19] = 16'hFFCE;
        rom[127][20] = 16'h0002;
        rom[127][21] = 16'h0010;
        rom[127][22] = 16'h0008;
        rom[127][23] = 16'hFFE7;
        rom[127][24] = 16'h001A;
        rom[127][25] = 16'hFFF4;
        rom[127][26] = 16'hFFE9;
        rom[127][27] = 16'hFFE8;
        rom[127][28] = 16'h001A;
        rom[127][29] = 16'h000D;
        rom[127][30] = 16'hFFE4;
        rom[127][31] = 16'h0001;
        rom[127][32] = 16'hFFEF;
        rom[127][33] = 16'h0024;
        rom[127][34] = 16'hFFAB;
        rom[127][35] = 16'h000F;
        rom[127][36] = 16'hFFE6;
        rom[127][37] = 16'h0013;
        rom[127][38] = 16'hFFFA;
        rom[127][39] = 16'hFFFE;
        rom[127][40] = 16'h0009;
        rom[127][41] = 16'hFFD5;
        rom[127][42] = 16'h0006;
        rom[127][43] = 16'hFFD2;
        rom[127][44] = 16'hFFF6;
        rom[127][45] = 16'hFFD9;
        rom[127][46] = 16'hFFF0;
        rom[127][47] = 16'h0008;
        rom[127][48] = 16'hFFC8;
        rom[127][49] = 16'hFFFA;
        rom[127][50] = 16'hFFC8;
        rom[127][51] = 16'h0012;
        rom[127][52] = 16'hFFE3;
        rom[127][53] = 16'hFFE8;
        rom[127][54] = 16'hFFF3;
        rom[127][55] = 16'h0002;
        rom[127][56] = 16'hFFEB;
        rom[127][57] = 16'h000C;
        rom[127][58] = 16'h0005;
        rom[127][59] = 16'hFFE5;
        rom[127][60] = 16'h000F;
        rom[127][61] = 16'h002B;
        rom[127][62] = 16'hFFF7;
        rom[127][63] = 16'h0001;
        rom[127][64] = 16'h0015;
        rom[127][65] = 16'h0007;
        rom[127][66] = 16'hFFDD;
        rom[127][67] = 16'hFFFC;
        rom[127][68] = 16'hFFF9;
        rom[127][69] = 16'h0002;
        rom[127][70] = 16'h0007;
        rom[127][71] = 16'hFFE8;
        rom[127][72] = 16'h0000;
        rom[127][73] = 16'h000C;
        rom[127][74] = 16'h0011;
        rom[127][75] = 16'hFFF4;
        rom[127][76] = 16'hFFCC;
        rom[127][77] = 16'hFFEC;
        rom[127][78] = 16'hFFF9;
        rom[127][79] = 16'hFFEF;
        rom[127][80] = 16'hFFF9;
        rom[127][81] = 16'hFFF9;
        rom[127][82] = 16'hFFD7;
        rom[127][83] = 16'h0008;
        rom[127][84] = 16'h0002;
        rom[127][85] = 16'hFFE7;
        rom[127][86] = 16'h0011;
        rom[127][87] = 16'hFFCE;
        rom[127][88] = 16'h0009;
        rom[127][89] = 16'hFFF1;
        rom[127][90] = 16'hFFF9;
        rom[127][91] = 16'hFFD7;
        rom[127][92] = 16'h000D;
        rom[127][93] = 16'h000E;
        rom[127][94] = 16'h0028;
        rom[127][95] = 16'h001B;
        rom[127][96] = 16'h0002;
        rom[127][97] = 16'h000B;
        rom[127][98] = 16'h0005;
        rom[127][99] = 16'hFFFF;
        rom[127][100] = 16'hFFE5;
        rom[127][101] = 16'hFFF0;
        rom[127][102] = 16'hFFFA;
        rom[127][103] = 16'hFFF1;
        rom[127][104] = 16'h0018;
        rom[127][105] = 16'h0006;
        rom[127][106] = 16'h001D;
        rom[127][107] = 16'hFFE0;
        rom[127][108] = 16'hFFE1;
        rom[127][109] = 16'h000F;
        rom[127][110] = 16'hFFFE;
        rom[127][111] = 16'hFFFD;
        rom[127][112] = 16'hFFE5;
        rom[127][113] = 16'hFFF5;
        rom[127][114] = 16'hFFFE;
        rom[127][115] = 16'hFFFE;
        rom[127][116] = 16'hFFF2;
        rom[127][117] = 16'hFFE7;
        rom[127][118] = 16'hFFF9;
        rom[127][119] = 16'hFFE5;
        rom[127][120] = 16'h0034;
        rom[127][121] = 16'hFFCC;
        rom[127][122] = 16'hFFD6;
        rom[127][123] = 16'h0006;
        rom[127][124] = 16'hFFA6;
        rom[127][125] = 16'h0025;
        rom[127][126] = 16'hFFF6;
        rom[127][127] = 16'hFFE8;
        rom[128][0] = 16'hFFF7;
        rom[128][1] = 16'h0024;
        rom[128][2] = 16'hFFEA;
        rom[128][3] = 16'hFFFA;
        rom[128][4] = 16'hFFF9;
        rom[128][5] = 16'h0010;
        rom[128][6] = 16'h000C;
        rom[128][7] = 16'h0025;
        rom[128][8] = 16'h0002;
        rom[128][9] = 16'h0011;
        rom[128][10] = 16'hFFCE;
        rom[128][11] = 16'hFFC3;
        rom[128][12] = 16'h0002;
        rom[128][13] = 16'h002E;
        rom[128][14] = 16'h0009;
        rom[128][15] = 16'h0010;
        rom[128][16] = 16'hFFF9;
        rom[128][17] = 16'h002F;
        rom[128][18] = 16'h0019;
        rom[128][19] = 16'hFFF8;
        rom[128][20] = 16'hFF9F;
        rom[128][21] = 16'h0005;
        rom[128][22] = 16'h0014;
        rom[128][23] = 16'hFFD9;
        rom[128][24] = 16'hFFC8;
        rom[128][25] = 16'h0002;
        rom[128][26] = 16'hFFFF;
        rom[128][27] = 16'hFFCD;
        rom[128][28] = 16'h0002;
        rom[128][29] = 16'h001B;
        rom[128][30] = 16'hFFD9;
        rom[128][31] = 16'hFFFA;
        rom[128][32] = 16'h0011;
        rom[128][33] = 16'h001D;
        rom[128][34] = 16'hFFDA;
        rom[128][35] = 16'h0011;
        rom[128][36] = 16'h0010;
        rom[128][37] = 16'hFFF0;
        rom[128][38] = 16'h000B;
        rom[128][39] = 16'hFFDD;
        rom[128][40] = 16'h0024;
        rom[128][41] = 16'h0005;
        rom[128][42] = 16'h0001;
        rom[128][43] = 16'hFFEC;
        rom[128][44] = 16'hFFEB;
        rom[128][45] = 16'h0016;
        rom[128][46] = 16'h000A;
        rom[128][47] = 16'h0012;
        rom[128][48] = 16'h0021;
        rom[128][49] = 16'h0044;
        rom[128][50] = 16'h0029;
        rom[128][51] = 16'hFFB3;
        rom[128][52] = 16'h0017;
        rom[128][53] = 16'h0003;
        rom[128][54] = 16'hFFEB;
        rom[128][55] = 16'hFFF4;
        rom[128][56] = 16'hFFD1;
        rom[128][57] = 16'hFFFB;
        rom[128][58] = 16'h0003;
        rom[128][59] = 16'hFFEA;
        rom[128][60] = 16'hFFE1;
        rom[128][61] = 16'hFFFE;
        rom[128][62] = 16'h0007;
        rom[128][63] = 16'h0018;
        rom[128][64] = 16'hFFDF;
        rom[128][65] = 16'h000C;
        rom[128][66] = 16'hFFD8;
        rom[128][67] = 16'h0016;
        rom[128][68] = 16'h001A;
        rom[128][69] = 16'h0007;
        rom[128][70] = 16'h0012;
        rom[128][71] = 16'h000B;
        rom[128][72] = 16'hFFCD;
        rom[128][73] = 16'h001D;
        rom[128][74] = 16'hFFF4;
        rom[128][75] = 16'hFFFE;
        rom[128][76] = 16'hFFEA;
        rom[128][77] = 16'hFFE1;
        rom[128][78] = 16'hFFE2;
        rom[128][79] = 16'h0010;
        rom[128][80] = 16'h000A;
        rom[128][81] = 16'hFFF9;
        rom[128][82] = 16'h001F;
        rom[128][83] = 16'hFFE6;
        rom[128][84] = 16'h0003;
        rom[128][85] = 16'h000E;
        rom[128][86] = 16'hFFF9;
        rom[128][87] = 16'hFFE6;
        rom[128][88] = 16'hFFE3;
        rom[128][89] = 16'h0005;
        rom[128][90] = 16'h0013;
        rom[128][91] = 16'h0040;
        rom[128][92] = 16'hFFE5;
        rom[128][93] = 16'hFFEE;
        rom[128][94] = 16'h0013;
        rom[128][95] = 16'hFFFF;
        rom[128][96] = 16'hFFF9;
        rom[128][97] = 16'hFFE5;
        rom[128][98] = 16'hFFFA;
        rom[128][99] = 16'hFFEA;
        rom[128][100] = 16'hFFC3;
        rom[128][101] = 16'hFFF4;
        rom[128][102] = 16'h000A;
        rom[128][103] = 16'hFFE5;
        rom[128][104] = 16'hFFF6;
        rom[128][105] = 16'hFFD2;
        rom[128][106] = 16'h0002;
        rom[128][107] = 16'hFFFB;
        rom[128][108] = 16'h0006;
        rom[128][109] = 16'h0030;
        rom[128][110] = 16'hFFFF;
        rom[128][111] = 16'hFFF3;
        rom[128][112] = 16'hFFCE;
        rom[128][113] = 16'hFFFE;
        rom[128][114] = 16'hFFF4;
        rom[128][115] = 16'hFFF6;
        rom[128][116] = 16'h0049;
        rom[128][117] = 16'h0023;
        rom[128][118] = 16'hFFE2;
        rom[128][119] = 16'h0007;
        rom[128][120] = 16'hFFF4;
        rom[128][121] = 16'hFFF0;
        rom[128][122] = 16'hFFB5;
        rom[128][123] = 16'h0007;
        rom[128][124] = 16'h001F;
        rom[128][125] = 16'hFFF0;
        rom[128][126] = 16'h0000;
        rom[128][127] = 16'hFFE1;
        rom[129][0] = 16'h0014;
        rom[129][1] = 16'hFFCF;
        rom[129][2] = 16'h0003;
        rom[129][3] = 16'hFFFD;
        rom[129][4] = 16'hFFC8;
        rom[129][5] = 16'hFFFB;
        rom[129][6] = 16'hFFE9;
        rom[129][7] = 16'hFFF3;
        rom[129][8] = 16'hFFC8;
        rom[129][9] = 16'h0012;
        rom[129][10] = 16'h0007;
        rom[129][11] = 16'h0002;
        rom[129][12] = 16'hFFEA;
        rom[129][13] = 16'hFFDC;
        rom[129][14] = 16'hFFEB;
        rom[129][15] = 16'h000C;
        rom[129][16] = 16'hFFE6;
        rom[129][17] = 16'hFFED;
        rom[129][18] = 16'h0035;
        rom[129][19] = 16'hFFE5;
        rom[129][20] = 16'h0023;
        rom[129][21] = 16'h0034;
        rom[129][22] = 16'hFFFC;
        rom[129][23] = 16'hFFFE;
        rom[129][24] = 16'h000B;
        rom[129][25] = 16'h002B;
        rom[129][26] = 16'hFFED;
        rom[129][27] = 16'h0001;
        rom[129][28] = 16'hFFDF;
        rom[129][29] = 16'hFFD7;
        rom[129][30] = 16'hFFD2;
        rom[129][31] = 16'hFFCD;
        rom[129][32] = 16'h0002;
        rom[129][33] = 16'h001B;
        rom[129][34] = 16'hFFEC;
        rom[129][35] = 16'hFFF2;
        rom[129][36] = 16'hFFED;
        rom[129][37] = 16'hFFE6;
        rom[129][38] = 16'hFFDD;
        rom[129][39] = 16'h0028;
        rom[129][40] = 16'hFFE1;
        rom[129][41] = 16'h0004;
        rom[129][42] = 16'hFFA1;
        rom[129][43] = 16'hFFFB;
        rom[129][44] = 16'hFFF5;
        rom[129][45] = 16'hFFF9;
        rom[129][46] = 16'hFFEF;
        rom[129][47] = 16'hFFFE;
        rom[129][48] = 16'hFFDD;
        rom[129][49] = 16'hFFE5;
        rom[129][50] = 16'hFFEB;
        rom[129][51] = 16'h0024;
        rom[129][52] = 16'h0002;
        rom[129][53] = 16'hFFFC;
        rom[129][54] = 16'hFFF0;
        rom[129][55] = 16'hFFF1;
        rom[129][56] = 16'hFFBB;
        rom[129][57] = 16'hFFF6;
        rom[129][58] = 16'hFFF3;
        rom[129][59] = 16'hFFE8;
        rom[129][60] = 16'hFFE1;
        rom[129][61] = 16'hFFCD;
        rom[129][62] = 16'hFFF3;
        rom[129][63] = 16'hFFD8;
        rom[129][64] = 16'h000A;
        rom[129][65] = 16'h0006;
        rom[129][66] = 16'hFFCA;
        rom[129][67] = 16'hFFC7;
        rom[129][68] = 16'hFFE5;
        rom[129][69] = 16'h0001;
        rom[129][70] = 16'h0005;
        rom[129][71] = 16'h0004;
        rom[129][72] = 16'h0003;
        rom[129][73] = 16'hFFAF;
        rom[129][74] = 16'hFFC5;
        rom[129][75] = 16'h000D;
        rom[129][76] = 16'h0013;
        rom[129][77] = 16'hFFB5;
        rom[129][78] = 16'h0011;
        rom[129][79] = 16'hFFD0;
        rom[129][80] = 16'h0013;
        rom[129][81] = 16'h000F;
        rom[129][82] = 16'hFFCD;
        rom[129][83] = 16'hFFDD;
        rom[129][84] = 16'h0007;
        rom[129][85] = 16'h0006;
        rom[129][86] = 16'h0008;
        rom[129][87] = 16'h000C;
        rom[129][88] = 16'h0023;
        rom[129][89] = 16'hFFF3;
        rom[129][90] = 16'hFFFA;
        rom[129][91] = 16'hFFFB;
        rom[129][92] = 16'hFFE1;
        rom[129][93] = 16'hFFE2;
        rom[129][94] = 16'hFFEE;
        rom[129][95] = 16'h0002;
        rom[129][96] = 16'h0026;
        rom[129][97] = 16'hFFC4;
        rom[129][98] = 16'hFFE4;
        rom[129][99] = 16'hFFEB;
        rom[129][100] = 16'h0010;
        rom[129][101] = 16'h000C;
        rom[129][102] = 16'h0003;
        rom[129][103] = 16'h0001;
        rom[129][104] = 16'hFFD4;
        rom[129][105] = 16'hFFD1;
        rom[129][106] = 16'hFFD2;
        rom[129][107] = 16'h0005;
        rom[129][108] = 16'h0029;
        rom[129][109] = 16'h0011;
        rom[129][110] = 16'hFFA2;
        rom[129][111] = 16'hFFF4;
        rom[129][112] = 16'hFFFC;
        rom[129][113] = 16'hFFE0;
        rom[129][114] = 16'hFFF9;
        rom[129][115] = 16'hFFF5;
        rom[129][116] = 16'h002C;
        rom[129][117] = 16'hFFF3;
        rom[129][118] = 16'hFFF9;
        rom[129][119] = 16'hFFD2;
        rom[129][120] = 16'h0009;
        rom[129][121] = 16'h0017;
        rom[129][122] = 16'hFFFD;
        rom[129][123] = 16'hFFFE;
        rom[129][124] = 16'hFFD1;
        rom[129][125] = 16'hFFE9;
        rom[129][126] = 16'h000B;
        rom[129][127] = 16'h0004;
        rom[130][0] = 16'hFFC8;
        rom[130][1] = 16'hFFFE;
        rom[130][2] = 16'hFFF6;
        rom[130][3] = 16'hFFFA;
        rom[130][4] = 16'h0007;
        rom[130][5] = 16'hFFFD;
        rom[130][6] = 16'h002C;
        rom[130][7] = 16'h001E;
        rom[130][8] = 16'hFFEE;
        rom[130][9] = 16'hFFE7;
        rom[130][10] = 16'hFFD3;
        rom[130][11] = 16'h0007;
        rom[130][12] = 16'hFFD2;
        rom[130][13] = 16'hFFEA;
        rom[130][14] = 16'hFFF9;
        rom[130][15] = 16'hFFE8;
        rom[130][16] = 16'h0033;
        rom[130][17] = 16'h0015;
        rom[130][18] = 16'h0024;
        rom[130][19] = 16'hFFB5;
        rom[130][20] = 16'h0022;
        rom[130][21] = 16'hFFF7;
        rom[130][22] = 16'hFFBB;
        rom[130][23] = 16'hFFF7;
        rom[130][24] = 16'h002E;
        rom[130][25] = 16'hFFED;
        rom[130][26] = 16'h0014;
        rom[130][27] = 16'h0009;
        rom[130][28] = 16'hFFEF;
        rom[130][29] = 16'hFFFA;
        rom[130][30] = 16'hFFCF;
        rom[130][31] = 16'hFFF4;
        rom[130][32] = 16'hFFD1;
        rom[130][33] = 16'h0007;
        rom[130][34] = 16'hFFF7;
        rom[130][35] = 16'hFFE8;
        rom[130][36] = 16'h0007;
        rom[130][37] = 16'hFFD7;
        rom[130][38] = 16'h0023;
        rom[130][39] = 16'hFFDB;
        rom[130][40] = 16'h001E;
        rom[130][41] = 16'hFF9D;
        rom[130][42] = 16'hFFE6;
        rom[130][43] = 16'hFFF4;
        rom[130][44] = 16'hFFFB;
        rom[130][45] = 16'h0013;
        rom[130][46] = 16'h0031;
        rom[130][47] = 16'hFFE9;
        rom[130][48] = 16'hFFF1;
        rom[130][49] = 16'hFFFF;
        rom[130][50] = 16'h000C;
        rom[130][51] = 16'h0007;
        rom[130][52] = 16'h000D;
        rom[130][53] = 16'h0028;
        rom[130][54] = 16'h0011;
        rom[130][55] = 16'hFFEE;
        rom[130][56] = 16'hFFF5;
        rom[130][57] = 16'h0012;
        rom[130][58] = 16'h001F;
        rom[130][59] = 16'h001F;
        rom[130][60] = 16'hFFE9;
        rom[130][61] = 16'hFFDF;
        rom[130][62] = 16'h001B;
        rom[130][63] = 16'h0011;
        rom[130][64] = 16'hFFD2;
        rom[130][65] = 16'h001D;
        rom[130][66] = 16'h0007;
        rom[130][67] = 16'hFFD8;
        rom[130][68] = 16'h000C;
        rom[130][69] = 16'hFFD1;
        rom[130][70] = 16'h0002;
        rom[130][71] = 16'hFFF8;
        rom[130][72] = 16'hFFE3;
        rom[130][73] = 16'hFFDB;
        rom[130][74] = 16'h0013;
        rom[130][75] = 16'h0013;
        rom[130][76] = 16'h0017;
        rom[130][77] = 16'h0004;
        rom[130][78] = 16'hFFD7;
        rom[130][79] = 16'hFFFE;
        rom[130][80] = 16'h002C;
        rom[130][81] = 16'h0020;
        rom[130][82] = 16'h0007;
        rom[130][83] = 16'hFFCD;
        rom[130][84] = 16'hFFEF;
        rom[130][85] = 16'h0019;
        rom[130][86] = 16'hFFEF;
        rom[130][87] = 16'h0003;
        rom[130][88] = 16'hFFF9;
        rom[130][89] = 16'h0021;
        rom[130][90] = 16'h001F;
        rom[130][91] = 16'h002A;
        rom[130][92] = 16'h0016;
        rom[130][93] = 16'hFFD3;
        rom[130][94] = 16'h0021;
        rom[130][95] = 16'hFFC9;
        rom[130][96] = 16'hFFC8;
        rom[130][97] = 16'h0033;
        rom[130][98] = 16'hFFCC;
        rom[130][99] = 16'h000C;
        rom[130][100] = 16'hFFD9;
        rom[130][101] = 16'hFFA9;
        rom[130][102] = 16'h001D;
        rom[130][103] = 16'hFFDA;
        rom[130][104] = 16'hFFF7;
        rom[130][105] = 16'h0036;
        rom[130][106] = 16'h0020;
        rom[130][107] = 16'hFFE6;
        rom[130][108] = 16'hFFC3;
        rom[130][109] = 16'hFFBA;
        rom[130][110] = 16'hFFFC;
        rom[130][111] = 16'hFFCD;
        rom[130][112] = 16'h0004;
        rom[130][113] = 16'hFFFC;
        rom[130][114] = 16'hFFFA;
        rom[130][115] = 16'hFFF9;
        rom[130][116] = 16'hFFFD;
        rom[130][117] = 16'hFFDE;
        rom[130][118] = 16'h001E;
        rom[130][119] = 16'h001D;
        rom[130][120] = 16'hFFDD;
        rom[130][121] = 16'h000D;
        rom[130][122] = 16'h0011;
        rom[130][123] = 16'h0019;
        rom[130][124] = 16'h001B;
        rom[130][125] = 16'h0006;
        rom[130][126] = 16'h0010;
        rom[130][127] = 16'hFFEF;
        rom[131][0] = 16'hFFE3;
        rom[131][1] = 16'h001D;
        rom[131][2] = 16'hFFCC;
        rom[131][3] = 16'hFFF7;
        rom[131][4] = 16'hFFF3;
        rom[131][5] = 16'hFFDE;
        rom[131][6] = 16'h0024;
        rom[131][7] = 16'h0012;
        rom[131][8] = 16'hFFF9;
        rom[131][9] = 16'hFFE8;
        rom[131][10] = 16'hFFED;
        rom[131][11] = 16'h0024;
        rom[131][12] = 16'h0036;
        rom[131][13] = 16'hFFED;
        rom[131][14] = 16'hFFD2;
        rom[131][15] = 16'h001B;
        rom[131][16] = 16'h0012;
        rom[131][17] = 16'hFFD6;
        rom[131][18] = 16'hFFF4;
        rom[131][19] = 16'hFFDF;
        rom[131][20] = 16'hFFE7;
        rom[131][21] = 16'h0007;
        rom[131][22] = 16'hFFD0;
        rom[131][23] = 16'hFFEF;
        rom[131][24] = 16'hFFD2;
        rom[131][25] = 16'hFFFE;
        rom[131][26] = 16'hFFEB;
        rom[131][27] = 16'hFFFF;
        rom[131][28] = 16'h003C;
        rom[131][29] = 16'h0003;
        rom[131][30] = 16'h0002;
        rom[131][31] = 16'h0004;
        rom[131][32] = 16'hFFB6;
        rom[131][33] = 16'hFFB8;
        rom[131][34] = 16'h0014;
        rom[131][35] = 16'h0011;
        rom[131][36] = 16'h0025;
        rom[131][37] = 16'h000A;
        rom[131][38] = 16'hFFA8;
        rom[131][39] = 16'h0016;
        rom[131][40] = 16'h0004;
        rom[131][41] = 16'h000C;
        rom[131][42] = 16'hFFD4;
        rom[131][43] = 16'hFFD4;
        rom[131][44] = 16'hFFFE;
        rom[131][45] = 16'h0009;
        rom[131][46] = 16'hFFF9;
        rom[131][47] = 16'h0014;
        rom[131][48] = 16'h000A;
        rom[131][49] = 16'h0016;
        rom[131][50] = 16'hFFBA;
        rom[131][51] = 16'hFFB9;
        rom[131][52] = 16'hFFBC;
        rom[131][53] = 16'hFFC3;
        rom[131][54] = 16'h0006;
        rom[131][55] = 16'h002C;
        rom[131][56] = 16'h0008;
        rom[131][57] = 16'hFFEF;
        rom[131][58] = 16'h0007;
        rom[131][59] = 16'hFFE4;
        rom[131][60] = 16'h0024;
        rom[131][61] = 16'hFFEE;
        rom[131][62] = 16'h0024;
        rom[131][63] = 16'h000B;
        rom[131][64] = 16'h0018;
        rom[131][65] = 16'h0004;
        rom[131][66] = 16'hFFE1;
        rom[131][67] = 16'hFFD7;
        rom[131][68] = 16'hFFF9;
        rom[131][69] = 16'hFFF7;
        rom[131][70] = 16'hFFE1;
        rom[131][71] = 16'hFFC9;
        rom[131][72] = 16'h0010;
        rom[131][73] = 16'hFFF8;
        rom[131][74] = 16'h000F;
        rom[131][75] = 16'hFFBE;
        rom[131][76] = 16'h0019;
        rom[131][77] = 16'hFFD0;
        rom[131][78] = 16'h000B;
        rom[131][79] = 16'h000F;
        rom[131][80] = 16'h0016;
        rom[131][81] = 16'h0000;
        rom[131][82] = 16'hFFD9;
        rom[131][83] = 16'hFFFE;
        rom[131][84] = 16'hFFFE;
        rom[131][85] = 16'hFFD4;
        rom[131][86] = 16'h002F;
        rom[131][87] = 16'hFFAB;
        rom[131][88] = 16'hFFE0;
        rom[131][89] = 16'hFFFA;
        rom[131][90] = 16'hFFED;
        rom[131][91] = 16'hFFFB;
        rom[131][92] = 16'hFFE1;
        rom[131][93] = 16'h000C;
        rom[131][94] = 16'hFFD2;
        rom[131][95] = 16'h000C;
        rom[131][96] = 16'hFFF7;
        rom[131][97] = 16'hFFFD;
        rom[131][98] = 16'h0018;
        rom[131][99] = 16'h0014;
        rom[131][100] = 16'h0023;
        rom[131][101] = 16'h0000;
        rom[131][102] = 16'h0024;
        rom[131][103] = 16'hFFEA;
        rom[131][104] = 16'hFFC3;
        rom[131][105] = 16'hFFA2;
        rom[131][106] = 16'h0011;
        rom[131][107] = 16'h0011;
        rom[131][108] = 16'h0019;
        rom[131][109] = 16'h000A;
        rom[131][110] = 16'h000F;
        rom[131][111] = 16'h002D;
        rom[131][112] = 16'hFFDD;
        rom[131][113] = 16'h000C;
        rom[131][114] = 16'h000F;
        rom[131][115] = 16'h0038;
        rom[131][116] = 16'hFFEF;
        rom[131][117] = 16'h0016;
        rom[131][118] = 16'h001B;
        rom[131][119] = 16'h0024;
        rom[131][120] = 16'hFFC5;
        rom[131][121] = 16'h002D;
        rom[131][122] = 16'hFFFA;
        rom[131][123] = 16'hFFCA;
        rom[131][124] = 16'hFFF6;
        rom[131][125] = 16'hFFD5;
        rom[131][126] = 16'hFFCE;
        rom[131][127] = 16'hFFE1;
        rom[132][0] = 16'hFFD2;
        rom[132][1] = 16'h001B;
        rom[132][2] = 16'hFFED;
        rom[132][3] = 16'h0007;
        rom[132][4] = 16'hFFE9;
        rom[132][5] = 16'h001C;
        rom[132][6] = 16'h001C;
        rom[132][7] = 16'hFFF8;
        rom[132][8] = 16'hFFEE;
        rom[132][9] = 16'h0007;
        rom[132][10] = 16'h0017;
        rom[132][11] = 16'hFFE8;
        rom[132][12] = 16'hFFE1;
        rom[132][13] = 16'hFFBD;
        rom[132][14] = 16'h001C;
        rom[132][15] = 16'hFFD4;
        rom[132][16] = 16'h000A;
        rom[132][17] = 16'h0033;
        rom[132][18] = 16'hFFF4;
        rom[132][19] = 16'hFFD6;
        rom[132][20] = 16'hFFB0;
        rom[132][21] = 16'hFFE2;
        rom[132][22] = 16'h0002;
        rom[132][23] = 16'h0020;
        rom[132][24] = 16'hFFCD;
        rom[132][25] = 16'hFFE7;
        rom[132][26] = 16'hFFE1;
        rom[132][27] = 16'hFFF2;
        rom[132][28] = 16'h0004;
        rom[132][29] = 16'hFFEF;
        rom[132][30] = 16'h0023;
        rom[132][31] = 16'h0012;
        rom[132][32] = 16'hFFE6;
        rom[132][33] = 16'hFFED;
        rom[132][34] = 16'h0024;
        rom[132][35] = 16'hFFED;
        rom[132][36] = 16'hFFF4;
        rom[132][37] = 16'h0008;
        rom[132][38] = 16'hFFF7;
        rom[132][39] = 16'hFFF6;
        rom[132][40] = 16'hFFE5;
        rom[132][41] = 16'hFFAB;
        rom[132][42] = 16'h0016;
        rom[132][43] = 16'hFFE7;
        rom[132][44] = 16'hFFF5;
        rom[132][45] = 16'hFFE0;
        rom[132][46] = 16'h0017;
        rom[132][47] = 16'h0010;
        rom[132][48] = 16'hFFF1;
        rom[132][49] = 16'hFFF7;
        rom[132][50] = 16'hFFF4;
        rom[132][51] = 16'h000B;
        rom[132][52] = 16'hFFEA;
        rom[132][53] = 16'hFFFF;
        rom[132][54] = 16'h000C;
        rom[132][55] = 16'h002B;
        rom[132][56] = 16'h0001;
        rom[132][57] = 16'hFFDB;
        rom[132][58] = 16'h0009;
        rom[132][59] = 16'h002B;
        rom[132][60] = 16'hFFF9;
        rom[132][61] = 16'hFFEC;
        rom[132][62] = 16'h0003;
        rom[132][63] = 16'hFFFC;
        rom[132][64] = 16'hFFED;
        rom[132][65] = 16'hFFF1;
        rom[132][66] = 16'hFFDD;
        rom[132][67] = 16'hFFDD;
        rom[132][68] = 16'h000C;
        rom[132][69] = 16'hFFC8;
        rom[132][70] = 16'hFFF3;
        rom[132][71] = 16'hFFE6;
        rom[132][72] = 16'hFFD3;
        rom[132][73] = 16'hFFDA;
        rom[132][74] = 16'h000F;
        rom[132][75] = 16'hFFE2;
        rom[132][76] = 16'hFFC4;
        rom[132][77] = 16'h0024;
        rom[132][78] = 16'h0001;
        rom[132][79] = 16'hFFFB;
        rom[132][80] = 16'h001A;
        rom[132][81] = 16'hFFD4;
        rom[132][82] = 16'hFFFD;
        rom[132][83] = 16'hFFF7;
        rom[132][84] = 16'h0002;
        rom[132][85] = 16'h0026;
        rom[132][86] = 16'hFFE3;
        rom[132][87] = 16'hFFDD;
        rom[132][88] = 16'hFFBE;
        rom[132][89] = 16'h003E;
        rom[132][90] = 16'hFFFD;
        rom[132][91] = 16'h003B;
        rom[132][92] = 16'h000C;
        rom[132][93] = 16'hFFD5;
        rom[132][94] = 16'h000B;
        rom[132][95] = 16'h0016;
        rom[132][96] = 16'h0016;
        rom[132][97] = 16'hFFD7;
        rom[132][98] = 16'hFFCE;
        rom[132][99] = 16'hFFFB;
        rom[132][100] = 16'h0010;
        rom[132][101] = 16'hFFF3;
        rom[132][102] = 16'h0011;
        rom[132][103] = 16'hFFCE;
        rom[132][104] = 16'h0011;
        rom[132][105] = 16'h0038;
        rom[132][106] = 16'h000C;
        rom[132][107] = 16'hFFFC;
        rom[132][108] = 16'hFFDB;
        rom[132][109] = 16'hFFF6;
        rom[132][110] = 16'hFFE5;
        rom[132][111] = 16'hFFDC;
        rom[132][112] = 16'hFFA7;
        rom[132][113] = 16'hFFC6;
        rom[132][114] = 16'hFFE4;
        rom[132][115] = 16'hFFD4;
        rom[132][116] = 16'hFFCD;
        rom[132][117] = 16'h0008;
        rom[132][118] = 16'h0027;
        rom[132][119] = 16'hFFC6;
        rom[132][120] = 16'hFFE8;
        rom[132][121] = 16'hFFF8;
        rom[132][122] = 16'hFFE1;
        rom[132][123] = 16'h001C;
        rom[132][124] = 16'hFFFB;
        rom[132][125] = 16'hFFE9;
        rom[132][126] = 16'hFFF3;
        rom[132][127] = 16'hFFCE;
        rom[133][0] = 16'hFFE5;
        rom[133][1] = 16'hFFF8;
        rom[133][2] = 16'hFFFE;
        rom[133][3] = 16'h0024;
        rom[133][4] = 16'hFFE8;
        rom[133][5] = 16'hFFFD;
        rom[133][6] = 16'hFFC0;
        rom[133][7] = 16'hFFF4;
        rom[133][8] = 16'hFFC8;
        rom[133][9] = 16'hFFF6;
        rom[133][10] = 16'hFFC5;
        rom[133][11] = 16'hFFF9;
        rom[133][12] = 16'hFFD7;
        rom[133][13] = 16'h001A;
        rom[133][14] = 16'hFFFE;
        rom[133][15] = 16'h0002;
        rom[133][16] = 16'hFFEF;
        rom[133][17] = 16'h0002;
        rom[133][18] = 16'hFFE5;
        rom[133][19] = 16'h0020;
        rom[133][20] = 16'h0020;
        rom[133][21] = 16'hFFFE;
        rom[133][22] = 16'hFFF5;
        rom[133][23] = 16'hFFCE;
        rom[133][24] = 16'hFFF4;
        rom[133][25] = 16'h0002;
        rom[133][26] = 16'hFFFC;
        rom[133][27] = 16'h0012;
        rom[133][28] = 16'h0008;
        rom[133][29] = 16'hFFF3;
        rom[133][30] = 16'h0011;
        rom[133][31] = 16'hFFE1;
        rom[133][32] = 16'hFFF0;
        rom[133][33] = 16'hFFCB;
        rom[133][34] = 16'hFFFE;
        rom[133][35] = 16'h0007;
        rom[133][36] = 16'hFFDC;
        rom[133][37] = 16'hFFFE;
        rom[133][38] = 16'hFFF4;
        rom[133][39] = 16'h0001;
        rom[133][40] = 16'hFFD7;
        rom[133][41] = 16'hFFD2;
        rom[133][42] = 16'h0019;
        rom[133][43] = 16'hFFD6;
        rom[133][44] = 16'h001F;
        rom[133][45] = 16'hFFB1;
        rom[133][46] = 16'h0003;
        rom[133][47] = 16'h0005;
        rom[133][48] = 16'h0006;
        rom[133][49] = 16'hFFE8;
        rom[133][50] = 16'hFFEF;
        rom[133][51] = 16'hFFE7;
        rom[133][52] = 16'hFFB1;
        rom[133][53] = 16'hFFCE;
        rom[133][54] = 16'hFFDD;
        rom[133][55] = 16'hFFF5;
        rom[133][56] = 16'hFFFD;
        rom[133][57] = 16'hFFDC;
        rom[133][58] = 16'hFFCD;
        rom[133][59] = 16'h0024;
        rom[133][60] = 16'h0039;
        rom[133][61] = 16'h000F;
        rom[133][62] = 16'hFFFA;
        rom[133][63] = 16'hFFD7;
        rom[133][64] = 16'h000F;
        rom[133][65] = 16'h000C;
        rom[133][66] = 16'h0008;
        rom[133][67] = 16'h0000;
        rom[133][68] = 16'hFFF0;
        rom[133][69] = 16'h001A;
        rom[133][70] = 16'hFFEA;
        rom[133][71] = 16'hFFDB;
        rom[133][72] = 16'hFFE4;
        rom[133][73] = 16'hFFCC;
        rom[133][74] = 16'hFFEA;
        rom[133][75] = 16'hFFDA;
        rom[133][76] = 16'h000F;
        rom[133][77] = 16'h0011;
        rom[133][78] = 16'h0009;
        rom[133][79] = 16'hFFD3;
        rom[133][80] = 16'hFFF3;
        rom[133][81] = 16'hFFD1;
        rom[133][82] = 16'h0005;
        rom[133][83] = 16'hFFF5;
        rom[133][84] = 16'h000C;
        rom[133][85] = 16'h002C;
        rom[133][86] = 16'hFFF6;
        rom[133][87] = 16'hFFEA;
        rom[133][88] = 16'hFFFD;
        rom[133][89] = 16'hFFE3;
        rom[133][90] = 16'h0004;
        rom[133][91] = 16'hFFE5;
        rom[133][92] = 16'h000F;
        rom[133][93] = 16'hFFF6;
        rom[133][94] = 16'h0003;
        rom[133][95] = 16'h0007;
        rom[133][96] = 16'hFFDE;
        rom[133][97] = 16'hFFE0;
        rom[133][98] = 16'hFFE0;
        rom[133][99] = 16'hFFF9;
        rom[133][100] = 16'hFFEC;
        rom[133][101] = 16'hFFFE;
        rom[133][102] = 16'hFFE1;
        rom[133][103] = 16'hFFCB;
        rom[133][104] = 16'h0004;
        rom[133][105] = 16'hFFC4;
        rom[133][106] = 16'h0004;
        rom[133][107] = 16'hFFBC;
        rom[133][108] = 16'hFFCF;
        rom[133][109] = 16'h002E;
        rom[133][110] = 16'h0002;
        rom[133][111] = 16'h0001;
        rom[133][112] = 16'h000D;
        rom[133][113] = 16'h0000;
        rom[133][114] = 16'h0001;
        rom[133][115] = 16'hFFE8;
        rom[133][116] = 16'h0007;
        rom[133][117] = 16'h000A;
        rom[133][118] = 16'hFFC9;
        rom[133][119] = 16'hFFEF;
        rom[133][120] = 16'hFFE6;
        rom[133][121] = 16'hFFEA;
        rom[133][122] = 16'hFFCF;
        rom[133][123] = 16'h001F;
        rom[133][124] = 16'hFFE5;
        rom[133][125] = 16'hFFFB;
        rom[133][126] = 16'h0007;
        rom[133][127] = 16'hFFD2;
        rom[134][0] = 16'h0005;
        rom[134][1] = 16'h0013;
        rom[134][2] = 16'h0009;
        rom[134][3] = 16'h0003;
        rom[134][4] = 16'hFFCC;
        rom[134][5] = 16'hFFE4;
        rom[134][6] = 16'h0002;
        rom[134][7] = 16'h000B;
        rom[134][8] = 16'hFFDF;
        rom[134][9] = 16'h001B;
        rom[134][10] = 16'h001F;
        rom[134][11] = 16'hFFC3;
        rom[134][12] = 16'h000E;
        rom[134][13] = 16'h001A;
        rom[134][14] = 16'hFFE3;
        rom[134][15] = 16'h0005;
        rom[134][16] = 16'hFFB1;
        rom[134][17] = 16'h0012;
        rom[134][18] = 16'hFFE1;
        rom[134][19] = 16'h001E;
        rom[134][20] = 16'hFFEA;
        rom[134][21] = 16'h0011;
        rom[134][22] = 16'hFFF5;
        rom[134][23] = 16'h000E;
        rom[134][24] = 16'h0021;
        rom[134][25] = 16'hFFD7;
        rom[134][26] = 16'hFFE9;
        rom[134][27] = 16'hFFAF;
        rom[134][28] = 16'h001F;
        rom[134][29] = 16'h0012;
        rom[134][30] = 16'hFFFE;
        rom[134][31] = 16'h001F;
        rom[134][32] = 16'h000E;
        rom[134][33] = 16'h0009;
        rom[134][34] = 16'hFFEF;
        rom[134][35] = 16'h0018;
        rom[134][36] = 16'h000C;
        rom[134][37] = 16'hFFFA;
        rom[134][38] = 16'h0017;
        rom[134][39] = 16'h003D;
        rom[134][40] = 16'hFFFC;
        rom[134][41] = 16'h001C;
        rom[134][42] = 16'h0006;
        rom[134][43] = 16'hFFDC;
        rom[134][44] = 16'hFFE2;
        rom[134][45] = 16'hFFFB;
        rom[134][46] = 16'hFFE1;
        rom[134][47] = 16'h0000;
        rom[134][48] = 16'hFFFE;
        rom[134][49] = 16'h0024;
        rom[134][50] = 16'h0031;
        rom[134][51] = 16'hFFF0;
        rom[134][52] = 16'h0011;
        rom[134][53] = 16'hFFFF;
        rom[134][54] = 16'hFFD8;
        rom[134][55] = 16'hFFCA;
        rom[134][56] = 16'h0006;
        rom[134][57] = 16'h0011;
        rom[134][58] = 16'hFFE1;
        rom[134][59] = 16'hFFC5;
        rom[134][60] = 16'hFFCC;
        rom[134][61] = 16'hFFF7;
        rom[134][62] = 16'hFFDF;
        rom[134][63] = 16'h0006;
        rom[134][64] = 16'hFFDE;
        rom[134][65] = 16'h0011;
        rom[134][66] = 16'hFFF4;
        rom[134][67] = 16'hFFEC;
        rom[134][68] = 16'hFFF6;
        rom[134][69] = 16'hFFE2;
        rom[134][70] = 16'h0020;
        rom[134][71] = 16'hFFC9;
        rom[134][72] = 16'h0016;
        rom[134][73] = 16'hFFF0;
        rom[134][74] = 16'h0015;
        rom[134][75] = 16'h0016;
        rom[134][76] = 16'h0024;
        rom[134][77] = 16'hFFE7;
        rom[134][78] = 16'hFFEF;
        rom[134][79] = 16'hFFAB;
        rom[134][80] = 16'hFFFA;
        rom[134][81] = 16'h0007;
        rom[134][82] = 16'hFFF7;
        rom[134][83] = 16'h0014;
        rom[134][84] = 16'h0012;
        rom[134][85] = 16'hFFEC;
        rom[134][86] = 16'h0010;
        rom[134][87] = 16'hFFCC;
        rom[134][88] = 16'hFFF0;
        rom[134][89] = 16'hFFD5;
        rom[134][90] = 16'h0000;
        rom[134][91] = 16'hFFA1;
        rom[134][92] = 16'hFFE5;
        rom[134][93] = 16'hFFFF;
        rom[134][94] = 16'h002B;
        rom[134][95] = 16'hFFDF;
        rom[134][96] = 16'hFFD9;
        rom[134][97] = 16'hFFDA;
        rom[134][98] = 16'hFFD7;
        rom[134][99] = 16'hFFEA;
        rom[134][100] = 16'hFFED;
        rom[134][101] = 16'hFFFF;
        rom[134][102] = 16'hFFF9;
        rom[134][103] = 16'hFFE5;
        rom[134][104] = 16'hFFD3;
        rom[134][105] = 16'hFFDE;
        rom[134][106] = 16'h0014;
        rom[134][107] = 16'hFFE4;
        rom[134][108] = 16'hFFEF;
        rom[134][109] = 16'hFFE9;
        rom[134][110] = 16'hFFF3;
        rom[134][111] = 16'h0004;
        rom[134][112] = 16'h0002;
        rom[134][113] = 16'h000C;
        rom[134][114] = 16'hFFFE;
        rom[134][115] = 16'hFFE9;
        rom[134][116] = 16'hFFD8;
        rom[134][117] = 16'h0007;
        rom[134][118] = 16'h000C;
        rom[134][119] = 16'hFFFD;
        rom[134][120] = 16'hFFF7;
        rom[134][121] = 16'h0002;
        rom[134][122] = 16'hFFCD;
        rom[134][123] = 16'hFFEC;
        rom[134][124] = 16'hFFF3;
        rom[134][125] = 16'hFFCD;
        rom[134][126] = 16'hFFD3;
        rom[134][127] = 16'hFFEF;
        rom[135][0] = 16'hFFF7;
        rom[135][1] = 16'h0013;
        rom[135][2] = 16'hFFD6;
        rom[135][3] = 16'hFFEF;
        rom[135][4] = 16'h0031;
        rom[135][5] = 16'h0012;
        rom[135][6] = 16'hFFF6;
        rom[135][7] = 16'h0002;
        rom[135][8] = 16'h0018;
        rom[135][9] = 16'hFFFD;
        rom[135][10] = 16'h0007;
        rom[135][11] = 16'hFF97;
        rom[135][12] = 16'h0010;
        rom[135][13] = 16'h001E;
        rom[135][14] = 16'h0002;
        rom[135][15] = 16'hFFFF;
        rom[135][16] = 16'hFFF1;
        rom[135][17] = 16'hFFF9;
        rom[135][18] = 16'hFFF4;
        rom[135][19] = 16'h0000;
        rom[135][20] = 16'h0006;
        rom[135][21] = 16'hFFE5;
        rom[135][22] = 16'hFFE2;
        rom[135][23] = 16'hFFF2;
        rom[135][24] = 16'hFFEC;
        rom[135][25] = 16'hFFF8;
        rom[135][26] = 16'hFFF0;
        rom[135][27] = 16'hFFE0;
        rom[135][28] = 16'hFFD2;
        rom[135][29] = 16'h0003;
        rom[135][30] = 16'h000C;
        rom[135][31] = 16'h0014;
        rom[135][32] = 16'hFFE1;
        rom[135][33] = 16'hFFDE;
        rom[135][34] = 16'hFFF4;
        rom[135][35] = 16'hFFF8;
        rom[135][36] = 16'h0017;
        rom[135][37] = 16'hFFDE;
        rom[135][38] = 16'hFFEA;
        rom[135][39] = 16'h0016;
        rom[135][40] = 16'h0021;
        rom[135][41] = 16'h0022;
        rom[135][42] = 16'h000B;
        rom[135][43] = 16'hFFE2;
        rom[135][44] = 16'h001B;
        rom[135][45] = 16'hFFD5;
        rom[135][46] = 16'h0009;
        rom[135][47] = 16'hFFEF;
        rom[135][48] = 16'h0010;
        rom[135][49] = 16'h0017;
        rom[135][50] = 16'hFFEF;
        rom[135][51] = 16'h0002;
        rom[135][52] = 16'hFFBF;
        rom[135][53] = 16'h000C;
        rom[135][54] = 16'h0002;
        rom[135][55] = 16'h0015;
        rom[135][56] = 16'h0011;
        rom[135][57] = 16'h001A;
        rom[135][58] = 16'h000E;
        rom[135][59] = 16'hFFDF;
        rom[135][60] = 16'hFFF9;
        rom[135][61] = 16'h0016;
        rom[135][62] = 16'h000C;
        rom[135][63] = 16'h0002;
        rom[135][64] = 16'hFFD6;
        rom[135][65] = 16'h0017;
        rom[135][66] = 16'hFFFB;
        rom[135][67] = 16'h0013;
        rom[135][68] = 16'hFFF8;
        rom[135][69] = 16'h0018;
        rom[135][70] = 16'hFFE3;
        rom[135][71] = 16'hFFBC;
        rom[135][72] = 16'hFFC7;
        rom[135][73] = 16'h0022;
        rom[135][74] = 16'h0007;
        rom[135][75] = 16'hFFE8;
        rom[135][76] = 16'hFFA1;
        rom[135][77] = 16'h0019;
        rom[135][78] = 16'h0006;
        rom[135][79] = 16'h0020;
        rom[135][80] = 16'h0020;
        rom[135][81] = 16'hFFEE;
        rom[135][82] = 16'h0013;
        rom[135][83] = 16'h0037;
        rom[135][84] = 16'hFFCD;
        rom[135][85] = 16'h0014;
        rom[135][86] = 16'h0007;
        rom[135][87] = 16'h0006;
        rom[135][88] = 16'h0007;
        rom[135][89] = 16'h0018;
        rom[135][90] = 16'hFFF6;
        rom[135][91] = 16'hFFEA;
        rom[135][92] = 16'hFFD9;
        rom[135][93] = 16'h0005;
        rom[135][94] = 16'h0018;
        rom[135][95] = 16'hFFFA;
        rom[135][96] = 16'hFFFE;
        rom[135][97] = 16'hFFFE;
        rom[135][98] = 16'h0024;
        rom[135][99] = 16'hFFF0;
        rom[135][100] = 16'hFFDC;
        rom[135][101] = 16'hFFDC;
        rom[135][102] = 16'h000C;
        rom[135][103] = 16'hFFF3;
        rom[135][104] = 16'h001E;
        rom[135][105] = 16'h0018;
        rom[135][106] = 16'hFFF1;
        rom[135][107] = 16'hFFF3;
        rom[135][108] = 16'hFFBA;
        rom[135][109] = 16'hFFBA;
        rom[135][110] = 16'h0009;
        rom[135][111] = 16'h0016;
        rom[135][112] = 16'h0016;
        rom[135][113] = 16'h001F;
        rom[135][114] = 16'hFFED;
        rom[135][115] = 16'hFFFE;
        rom[135][116] = 16'hFFF0;
        rom[135][117] = 16'h0006;
        rom[135][118] = 16'h0027;
        rom[135][119] = 16'hFFD3;
        rom[135][120] = 16'hFFCD;
        rom[135][121] = 16'h0016;
        rom[135][122] = 16'hFFE4;
        rom[135][123] = 16'hFFC3;
        rom[135][124] = 16'hFFD4;
        rom[135][125] = 16'hFFEE;
        rom[135][126] = 16'hFFEF;
        rom[135][127] = 16'h000D;
        rom[136][0] = 16'h0009;
        rom[136][1] = 16'h000C;
        rom[136][2] = 16'h001B;
        rom[136][3] = 16'hFFE8;
        rom[136][4] = 16'hFFF2;
        rom[136][5] = 16'hFFFE;
        rom[136][6] = 16'hFFF4;
        rom[136][7] = 16'h0037;
        rom[136][8] = 16'h001D;
        rom[136][9] = 16'hFFEA;
        rom[136][10] = 16'hFFD6;
        rom[136][11] = 16'hFFE0;
        rom[136][12] = 16'hFFE6;
        rom[136][13] = 16'hFFFA;
        rom[136][14] = 16'hFFEB;
        rom[136][15] = 16'h0028;
        rom[136][16] = 16'hFFB8;
        rom[136][17] = 16'h0015;
        rom[136][18] = 16'hFFEE;
        rom[136][19] = 16'h0016;
        rom[136][20] = 16'h000B;
        rom[136][21] = 16'h001B;
        rom[136][22] = 16'h0002;
        rom[136][23] = 16'h0005;
        rom[136][24] = 16'h0003;
        rom[136][25] = 16'hFFEC;
        rom[136][26] = 16'h0032;
        rom[136][27] = 16'hFFC0;
        rom[136][28] = 16'hFFE0;
        rom[136][29] = 16'hFFF8;
        rom[136][30] = 16'hFFF4;
        rom[136][31] = 16'h0012;
        rom[136][32] = 16'h0002;
        rom[136][33] = 16'h0006;
        rom[136][34] = 16'hFFEF;
        rom[136][35] = 16'hFFE2;
        rom[136][36] = 16'h0029;
        rom[136][37] = 16'h0007;
        rom[136][38] = 16'h0016;
        rom[136][39] = 16'hFFB5;
        rom[136][40] = 16'hFFDB;
        rom[136][41] = 16'h000F;
        rom[136][42] = 16'h000C;
        rom[136][43] = 16'hFFD4;
        rom[136][44] = 16'hFFE5;
        rom[136][45] = 16'hFFF8;
        rom[136][46] = 16'h0009;
        rom[136][47] = 16'hFFF7;
        rom[136][48] = 16'hFFEA;
        rom[136][49] = 16'h0032;
        rom[136][50] = 16'h0008;
        rom[136][51] = 16'hFFE0;
        rom[136][52] = 16'h002B;
        rom[136][53] = 16'h000C;
        rom[136][54] = 16'hFFF0;
        rom[136][55] = 16'h0011;
        rom[136][56] = 16'h0001;
        rom[136][57] = 16'hFFE0;
        rom[136][58] = 16'h000E;
        rom[136][59] = 16'hFFCC;
        rom[136][60] = 16'hFFF9;
        rom[136][61] = 16'h000F;
        rom[136][62] = 16'hFFD7;
        rom[136][63] = 16'h0019;
        rom[136][64] = 16'hFFF7;
        rom[136][65] = 16'h0018;
        rom[136][66] = 16'h0018;
        rom[136][67] = 16'hFFF4;
        rom[136][68] = 16'hFFE9;
        rom[136][69] = 16'h0002;
        rom[136][70] = 16'h001B;
        rom[136][71] = 16'hFFFB;
        rom[136][72] = 16'hFFF1;
        rom[136][73] = 16'hFFD5;
        rom[136][74] = 16'h0011;
        rom[136][75] = 16'h0004;
        rom[136][76] = 16'h000A;
        rom[136][77] = 16'hFFD1;
        rom[136][78] = 16'hFFEF;
        rom[136][79] = 16'hFFFD;
        rom[136][80] = 16'h002E;
        rom[136][81] = 16'hFFF1;
        rom[136][82] = 16'h000F;
        rom[136][83] = 16'hFFD9;
        rom[136][84] = 16'h0002;
        rom[136][85] = 16'hFFF3;
        rom[136][86] = 16'hFFDC;
        rom[136][87] = 16'hFFD7;
        rom[136][88] = 16'h000E;
        rom[136][89] = 16'hFFCF;
        rom[136][90] = 16'h0024;
        rom[136][91] = 16'hFFEA;
        rom[136][92] = 16'h0007;
        rom[136][93] = 16'h000C;
        rom[136][94] = 16'hFFF0;
        rom[136][95] = 16'h0004;
        rom[136][96] = 16'hFFC4;
        rom[136][97] = 16'hFFDA;
        rom[136][98] = 16'hFFDF;
        rom[136][99] = 16'h002C;
        rom[136][100] = 16'hFFA8;
        rom[136][101] = 16'hFFD9;
        rom[136][102] = 16'hFFFE;
        rom[136][103] = 16'hFFF5;
        rom[136][104] = 16'hFFEB;
        rom[136][105] = 16'hFFB7;
        rom[136][106] = 16'hFFF9;
        rom[136][107] = 16'hFFF0;
        rom[136][108] = 16'h0007;
        rom[136][109] = 16'h0004;
        rom[136][110] = 16'h0002;
        rom[136][111] = 16'h0024;
        rom[136][112] = 16'hFFBC;
        rom[136][113] = 16'hFFFE;
        rom[136][114] = 16'hFFEA;
        rom[136][115] = 16'hFFDB;
        rom[136][116] = 16'h0007;
        rom[136][117] = 16'h001B;
        rom[136][118] = 16'hFFE8;
        rom[136][119] = 16'hFFFF;
        rom[136][120] = 16'hFFCC;
        rom[136][121] = 16'hFFBB;
        rom[136][122] = 16'hFFC4;
        rom[136][123] = 16'hFFF8;
        rom[136][124] = 16'h0001;
        rom[136][125] = 16'hFFCE;
        rom[136][126] = 16'h0009;
        rom[136][127] = 16'hFFF8;
        rom[137][0] = 16'h003D;
        rom[137][1] = 16'hFFF6;
        rom[137][2] = 16'hFFD9;
        rom[137][3] = 16'hFFE5;
        rom[137][4] = 16'hFFD7;
        rom[137][5] = 16'h000C;
        rom[137][6] = 16'h0019;
        rom[137][7] = 16'hFFD6;
        rom[137][8] = 16'hFFE9;
        rom[137][9] = 16'hFFC4;
        rom[137][10] = 16'h0002;
        rom[137][11] = 16'hFFFA;
        rom[137][12] = 16'h0004;
        rom[137][13] = 16'hFFED;
        rom[137][14] = 16'hFFEA;
        rom[137][15] = 16'hFFDC;
        rom[137][16] = 16'hFFF6;
        rom[137][17] = 16'h0029;
        rom[137][18] = 16'hFFF0;
        rom[137][19] = 16'h0002;
        rom[137][20] = 16'hFFF4;
        rom[137][21] = 16'hFFD4;
        rom[137][22] = 16'h000D;
        rom[137][23] = 16'hFFCD;
        rom[137][24] = 16'h0066;
        rom[137][25] = 16'hFFA0;
        rom[137][26] = 16'h001D;
        rom[137][27] = 16'hFFBB;
        rom[137][28] = 16'h0025;
        rom[137][29] = 16'h0005;
        rom[137][30] = 16'hFFFE;
        rom[137][31] = 16'hFFDA;
        rom[137][32] = 16'h0022;
        rom[137][33] = 16'hFFC2;
        rom[137][34] = 16'h0003;
        rom[137][35] = 16'hFFFB;
        rom[137][36] = 16'h000C;
        rom[137][37] = 16'hFFEF;
        rom[137][38] = 16'hFFCD;
        rom[137][39] = 16'h0016;
        rom[137][40] = 16'hFFF4;
        rom[137][41] = 16'h0014;
        rom[137][42] = 16'hFFFE;
        rom[137][43] = 16'hFFEA;
        rom[137][44] = 16'hFFF1;
        rom[137][45] = 16'hFFEA;
        rom[137][46] = 16'h0011;
        rom[137][47] = 16'hFFCF;
        rom[137][48] = 16'h0011;
        rom[137][49] = 16'h0002;
        rom[137][50] = 16'hFFD5;
        rom[137][51] = 16'h0008;
        rom[137][52] = 16'h0014;
        rom[137][53] = 16'h0005;
        rom[137][54] = 16'h0006;
        rom[137][55] = 16'hFFF1;
        rom[137][56] = 16'h0002;
        rom[137][57] = 16'hFFFE;
        rom[137][58] = 16'hFFDA;
        rom[137][59] = 16'hFFE9;
        rom[137][60] = 16'h0008;
        rom[137][61] = 16'hFFD8;
        rom[137][62] = 16'hFFE7;
        rom[137][63] = 16'hFFE9;
        rom[137][64] = 16'h000F;
        rom[137][65] = 16'h0007;
        rom[137][66] = 16'h001F;
        rom[137][67] = 16'h000B;
        rom[137][68] = 16'h002B;
        rom[137][69] = 16'h0002;
        rom[137][70] = 16'h0004;
        rom[137][71] = 16'h0022;
        rom[137][72] = 16'hFFF4;
        rom[137][73] = 16'h000C;
        rom[137][74] = 16'h000C;
        rom[137][75] = 16'hFFCA;
        rom[137][76] = 16'h0068;
        rom[137][77] = 16'h001F;
        rom[137][78] = 16'h0007;
        rom[137][79] = 16'hFFEB;
        rom[137][80] = 16'h0000;
        rom[137][81] = 16'hFFFD;
        rom[137][82] = 16'hFFCB;
        rom[137][83] = 16'h0004;
        rom[137][84] = 16'hFFF9;
        rom[137][85] = 16'h0002;
        rom[137][86] = 16'h0013;
        rom[137][87] = 16'h0003;
        rom[137][88] = 16'h000B;
        rom[137][89] = 16'h0016;
        rom[137][90] = 16'hFFF4;
        rom[137][91] = 16'h0020;
        rom[137][92] = 16'hFF99;
        rom[137][93] = 16'h003D;
        rom[137][94] = 16'h0011;
        rom[137][95] = 16'h0043;
        rom[137][96] = 16'h0014;
        rom[137][97] = 16'h000F;
        rom[137][98] = 16'h0010;
        rom[137][99] = 16'h0024;
        rom[137][100] = 16'h0034;
        rom[137][101] = 16'h0030;
        rom[137][102] = 16'hFFE7;
        rom[137][103] = 16'h0014;
        rom[137][104] = 16'h002A;
        rom[137][105] = 16'hFFF9;
        rom[137][106] = 16'hFFEF;
        rom[137][107] = 16'h0016;
        rom[137][108] = 16'hFFD4;
        rom[137][109] = 16'h0012;
        rom[137][110] = 16'hFFF1;
        rom[137][111] = 16'h0014;
        rom[137][112] = 16'hFFF2;
        rom[137][113] = 16'hFFD3;
        rom[137][114] = 16'h0001;
        rom[137][115] = 16'hFFF7;
        rom[137][116] = 16'hFFBD;
        rom[137][117] = 16'h0012;
        rom[137][118] = 16'hFFED;
        rom[137][119] = 16'hFFE0;
        rom[137][120] = 16'h000A;
        rom[137][121] = 16'hFFE2;
        rom[137][122] = 16'hFFF4;
        rom[137][123] = 16'hFFC0;
        rom[137][124] = 16'h0023;
        rom[137][125] = 16'h000C;
        rom[137][126] = 16'h0014;
        rom[137][127] = 16'h000A;
        rom[138][0] = 16'hFFCD;
        rom[138][1] = 16'hFFFE;
        rom[138][2] = 16'h000B;
        rom[138][3] = 16'h0002;
        rom[138][4] = 16'h002D;
        rom[138][5] = 16'h0009;
        rom[138][6] = 16'hFFF1;
        rom[138][7] = 16'h0011;
        rom[138][8] = 16'h0029;
        rom[138][9] = 16'hFFE3;
        rom[138][10] = 16'hFFDC;
        rom[138][11] = 16'hFFF0;
        rom[138][12] = 16'hFFF4;
        rom[138][13] = 16'hFFDC;
        rom[138][14] = 16'hFFEF;
        rom[138][15] = 16'h0013;
        rom[138][16] = 16'h0004;
        rom[138][17] = 16'h0006;
        rom[138][18] = 16'h0015;
        rom[138][19] = 16'h002B;
        rom[138][20] = 16'hFFF9;
        rom[138][21] = 16'hFFD4;
        rom[138][22] = 16'hFFEC;
        rom[138][23] = 16'h000C;
        rom[138][24] = 16'hFFCA;
        rom[138][25] = 16'h0016;
        rom[138][26] = 16'h0003;
        rom[138][27] = 16'hFFD5;
        rom[138][28] = 16'h0028;
        rom[138][29] = 16'h000E;
        rom[138][30] = 16'hFFF6;
        rom[138][31] = 16'hFFB8;
        rom[138][32] = 16'h0010;
        rom[138][33] = 16'hFFE5;
        rom[138][34] = 16'hFFDD;
        rom[138][35] = 16'hFFF1;
        rom[138][36] = 16'h0014;
        rom[138][37] = 16'h0002;
        rom[138][38] = 16'hFFCC;
        rom[138][39] = 16'hFFE3;
        rom[138][40] = 16'hFFFC;
        rom[138][41] = 16'hFFF8;
        rom[138][42] = 16'hFFDD;
        rom[138][43] = 16'h0003;
        rom[138][44] = 16'hFFE5;
        rom[138][45] = 16'h000C;
        rom[138][46] = 16'h001F;
        rom[138][47] = 16'h0040;
        rom[138][48] = 16'h000A;
        rom[138][49] = 16'h003A;
        rom[138][50] = 16'hFFFB;
        rom[138][51] = 16'hFFE2;
        rom[138][52] = 16'hFFFB;
        rom[138][53] = 16'h0016;
        rom[138][54] = 16'hFFEB;
        rom[138][55] = 16'h001B;
        rom[138][56] = 16'hFFEE;
        rom[138][57] = 16'hFFDE;
        rom[138][58] = 16'hFFFC;
        rom[138][59] = 16'h0035;
        rom[138][60] = 16'h0011;
        rom[138][61] = 16'hFFD0;
        rom[138][62] = 16'h0033;
        rom[138][63] = 16'hFFFE;
        rom[138][64] = 16'h0007;
        rom[138][65] = 16'hFFF3;
        rom[138][66] = 16'hFFF7;
        rom[138][67] = 16'hFFE4;
        rom[138][68] = 16'hFFE4;
        rom[138][69] = 16'h000C;
        rom[138][70] = 16'hFFD0;
        rom[138][71] = 16'hFFF2;
        rom[138][72] = 16'hFFFE;
        rom[138][73] = 16'hFFF3;
        rom[138][74] = 16'hFFCA;
        rom[138][75] = 16'hFFEA;
        rom[138][76] = 16'h0018;
        rom[138][77] = 16'hFFEF;
        rom[138][78] = 16'hFFF4;
        rom[138][79] = 16'h000B;
        rom[138][80] = 16'h0002;
        rom[138][81] = 16'h0023;
        rom[138][82] = 16'h0016;
        rom[138][83] = 16'h002D;
        rom[138][84] = 16'h0019;
        rom[138][85] = 16'hFFF9;
        rom[138][86] = 16'hFFD3;
        rom[138][87] = 16'hFFDC;
        rom[138][88] = 16'h0016;
        rom[138][89] = 16'h001B;
        rom[138][90] = 16'h001B;
        rom[138][91] = 16'hFFDA;
        rom[138][92] = 16'hFFED;
        rom[138][93] = 16'hFFD9;
        rom[138][94] = 16'hFFFB;
        rom[138][95] = 16'hFFF9;
        rom[138][96] = 16'hFFEC;
        rom[138][97] = 16'hFFF4;
        rom[138][98] = 16'hFFF9;
        rom[138][99] = 16'h000C;
        rom[138][100] = 16'hFFF1;
        rom[138][101] = 16'hFFEF;
        rom[138][102] = 16'hFFED;
        rom[138][103] = 16'hFFFE;
        rom[138][104] = 16'hFFEB;
        rom[138][105] = 16'hFFDA;
        rom[138][106] = 16'h000D;
        rom[138][107] = 16'h001B;
        rom[138][108] = 16'hFFDD;
        rom[138][109] = 16'hFFFA;
        rom[138][110] = 16'h0022;
        rom[138][111] = 16'h0031;
        rom[138][112] = 16'hFFF5;
        rom[138][113] = 16'hFFFE;
        rom[138][114] = 16'hFFEA;
        rom[138][115] = 16'h000E;
        rom[138][116] = 16'h0002;
        rom[138][117] = 16'h0005;
        rom[138][118] = 16'h0011;
        rom[138][119] = 16'h0008;
        rom[138][120] = 16'hFFDA;
        rom[138][121] = 16'hFFF9;
        rom[138][122] = 16'hFFFF;
        rom[138][123] = 16'h0017;
        rom[138][124] = 16'hFFF3;
        rom[138][125] = 16'hFFFD;
        rom[138][126] = 16'hFFD2;
        rom[138][127] = 16'hFFF1;
        rom[139][0] = 16'h0016;
        rom[139][1] = 16'hFFF7;
        rom[139][2] = 16'hFFC8;
        rom[139][3] = 16'hFFFD;
        rom[139][4] = 16'h0030;
        rom[139][5] = 16'h001F;
        rom[139][6] = 16'hFFD2;
        rom[139][7] = 16'h0016;
        rom[139][8] = 16'h001D;
        rom[139][9] = 16'h000D;
        rom[139][10] = 16'hFFC6;
        rom[139][11] = 16'hFFC3;
        rom[139][12] = 16'hFFD8;
        rom[139][13] = 16'h001F;
        rom[139][14] = 16'hFFEC;
        rom[139][15] = 16'h002A;
        rom[139][16] = 16'hFFCC;
        rom[139][17] = 16'hFFF4;
        rom[139][18] = 16'h0000;
        rom[139][19] = 16'h0011;
        rom[139][20] = 16'h0031;
        rom[139][21] = 16'hFFF8;
        rom[139][22] = 16'hFFF0;
        rom[139][23] = 16'hFFFE;
        rom[139][24] = 16'h001B;
        rom[139][25] = 16'hFFF6;
        rom[139][26] = 16'hFFE6;
        rom[139][27] = 16'h0008;
        rom[139][28] = 16'h0016;
        rom[139][29] = 16'h0016;
        rom[139][30] = 16'h0027;
        rom[139][31] = 16'h000C;
        rom[139][32] = 16'hFFD9;
        rom[139][33] = 16'hFFE5;
        rom[139][34] = 16'hFFF0;
        rom[139][35] = 16'h000C;
        rom[139][36] = 16'hFFF5;
        rom[139][37] = 16'hFFF7;
        rom[139][38] = 16'h001F;
        rom[139][39] = 16'hFFFB;
        rom[139][40] = 16'hFFDC;
        rom[139][41] = 16'h000A;
        rom[139][42] = 16'hFFE8;
        rom[139][43] = 16'hFFC3;
        rom[139][44] = 16'hFFF5;
        rom[139][45] = 16'hFFF5;
        rom[139][46] = 16'hFFEB;
        rom[139][47] = 16'hFFFF;
        rom[139][48] = 16'hFFEE;
        rom[139][49] = 16'hFFD6;
        rom[139][50] = 16'hFFF4;
        rom[139][51] = 16'h0016;
        rom[139][52] = 16'hFFD5;
        rom[139][53] = 16'hFFE9;
        rom[139][54] = 16'h0007;
        rom[139][55] = 16'hFFE2;
        rom[139][56] = 16'hFFE5;
        rom[139][57] = 16'hFFFF;
        rom[139][58] = 16'hFF9E;
        rom[139][59] = 16'h0015;
        rom[139][60] = 16'h001F;
        rom[139][61] = 16'h0001;
        rom[139][62] = 16'hFFF4;
        rom[139][63] = 16'h0007;
        rom[139][64] = 16'h0001;
        rom[139][65] = 16'hFFFD;
        rom[139][66] = 16'hFFFF;
        rom[139][67] = 16'h003B;
        rom[139][68] = 16'hFFFC;
        rom[139][69] = 16'hFFF2;
        rom[139][70] = 16'hFFE9;
        rom[139][71] = 16'hFFD0;
        rom[139][72] = 16'h0033;
        rom[139][73] = 16'hFFF8;
        rom[139][74] = 16'h0001;
        rom[139][75] = 16'hFFF6;
        rom[139][76] = 16'hFFF1;
        rom[139][77] = 16'hFFA3;
        rom[139][78] = 16'h000E;
        rom[139][79] = 16'hFFBF;
        rom[139][80] = 16'h002B;
        rom[139][81] = 16'hFFF0;
        rom[139][82] = 16'h0018;
        rom[139][83] = 16'h0015;
        rom[139][84] = 16'hFFD9;
        rom[139][85] = 16'hFFE7;
        rom[139][86] = 16'hFFEE;
        rom[139][87] = 16'hFFFB;
        rom[139][88] = 16'h001F;
        rom[139][89] = 16'hFFE7;
        rom[139][90] = 16'h0004;
        rom[139][91] = 16'hFFD5;
        rom[139][92] = 16'h0003;
        rom[139][93] = 16'h0007;
        rom[139][94] = 16'h0001;
        rom[139][95] = 16'h0006;
        rom[139][96] = 16'hFFE3;
        rom[139][97] = 16'hFFE8;
        rom[139][98] = 16'hFFE6;
        rom[139][99] = 16'h0020;
        rom[139][100] = 16'hFFD7;
        rom[139][101] = 16'hFFD7;
        rom[139][102] = 16'hFFDC;
        rom[139][103] = 16'h0017;
        rom[139][104] = 16'hFFEE;
        rom[139][105] = 16'h0015;
        rom[139][106] = 16'hFFD6;
        rom[139][107] = 16'h0004;
        rom[139][108] = 16'hFFCE;
        rom[139][109] = 16'h000D;
        rom[139][110] = 16'h0002;
        rom[139][111] = 16'hFFF5;
        rom[139][112] = 16'hFFE2;
        rom[139][113] = 16'hFFE4;
        rom[139][114] = 16'hFFF9;
        rom[139][115] = 16'hFFDC;
        rom[139][116] = 16'hFFE1;
        rom[139][117] = 16'h0006;
        rom[139][118] = 16'h0012;
        rom[139][119] = 16'h0003;
        rom[139][120] = 16'h0033;
        rom[139][121] = 16'hFFEE;
        rom[139][122] = 16'hFFC9;
        rom[139][123] = 16'h0008;
        rom[139][124] = 16'hFFE7;
        rom[139][125] = 16'h0010;
        rom[139][126] = 16'hFFDE;
        rom[139][127] = 16'hFFCC;
        rom[140][0] = 16'h0044;
        rom[140][1] = 16'hFFFD;
        rom[140][2] = 16'hFFC9;
        rom[140][3] = 16'hFFF9;
        rom[140][4] = 16'h001A;
        rom[140][5] = 16'hFFDC;
        rom[140][6] = 16'h0006;
        rom[140][7] = 16'h0000;
        rom[140][8] = 16'h0020;
        rom[140][9] = 16'hFFFF;
        rom[140][10] = 16'h0001;
        rom[140][11] = 16'h000C;
        rom[140][12] = 16'h0020;
        rom[140][13] = 16'h000F;
        rom[140][14] = 16'h0000;
        rom[140][15] = 16'h000E;
        rom[140][16] = 16'h0000;
        rom[140][17] = 16'hFFF9;
        rom[140][18] = 16'hFFF4;
        rom[140][19] = 16'hFFBD;
        rom[140][20] = 16'hFFF4;
        rom[140][21] = 16'h0014;
        rom[140][22] = 16'h0017;
        rom[140][23] = 16'h0011;
        rom[140][24] = 16'h0029;
        rom[140][25] = 16'hFFE8;
        rom[140][26] = 16'h0011;
        rom[140][27] = 16'hFFBE;
        rom[140][28] = 16'h0032;
        rom[140][29] = 16'hFFDD;
        rom[140][30] = 16'h001B;
        rom[140][31] = 16'hFFE1;
        rom[140][32] = 16'hFFC8;
        rom[140][33] = 16'hFFFB;
        rom[140][34] = 16'hFFF6;
        rom[140][35] = 16'hFFF4;
        rom[140][36] = 16'hFFF1;
        rom[140][37] = 16'hFFFE;
        rom[140][38] = 16'hFFFE;
        rom[140][39] = 16'h000F;
        rom[140][40] = 16'hFFCF;
        rom[140][41] = 16'hFFFC;
        rom[140][42] = 16'h0004;
        rom[140][43] = 16'hFF9E;
        rom[140][44] = 16'h0002;
        rom[140][45] = 16'hFFD1;
        rom[140][46] = 16'h0003;
        rom[140][47] = 16'hFFD0;
        rom[140][48] = 16'hFFE5;
        rom[140][49] = 16'hFFFA;
        rom[140][50] = 16'hFFD4;
        rom[140][51] = 16'h0009;
        rom[140][52] = 16'h000E;
        rom[140][53] = 16'hFFC8;
        rom[140][54] = 16'hFFD7;
        rom[140][55] = 16'hFFE2;
        rom[140][56] = 16'hFFE9;
        rom[140][57] = 16'h001D;
        rom[140][58] = 16'hFFE4;
        rom[140][59] = 16'hFFD5;
        rom[140][60] = 16'hFFFC;
        rom[140][61] = 16'hFFD1;
        rom[140][62] = 16'hFFFE;
        rom[140][63] = 16'hFFE9;
        rom[140][64] = 16'hFFEF;
        rom[140][65] = 16'h0021;
        rom[140][66] = 16'h0002;
        rom[140][67] = 16'h0002;
        rom[140][68] = 16'h0005;
        rom[140][69] = 16'hFFF9;
        rom[140][70] = 16'h0020;
        rom[140][71] = 16'h0004;
        rom[140][72] = 16'h000F;
        rom[140][73] = 16'hFFF2;
        rom[140][74] = 16'h0007;
        rom[140][75] = 16'h0013;
        rom[140][76] = 16'h000B;
        rom[140][77] = 16'hFFFD;
        rom[140][78] = 16'h0038;
        rom[140][79] = 16'h0001;
        rom[140][80] = 16'hFFF8;
        rom[140][81] = 16'hFFC3;
        rom[140][82] = 16'hFFE1;
        rom[140][83] = 16'hFFEB;
        rom[140][84] = 16'h0002;
        rom[140][85] = 16'hFFB8;
        rom[140][86] = 16'hFFD6;
        rom[140][87] = 16'h003D;
        rom[140][88] = 16'hFFE0;
        rom[140][89] = 16'h0010;
        rom[140][90] = 16'hFFE6;
        rom[140][91] = 16'h0030;
        rom[140][92] = 16'h002E;
        rom[140][93] = 16'h0020;
        rom[140][94] = 16'h001F;
        rom[140][95] = 16'h0019;
        rom[140][96] = 16'h002A;
        rom[140][97] = 16'h0023;
        rom[140][98] = 16'hFFE6;
        rom[140][99] = 16'h000B;
        rom[140][100] = 16'h0024;
        rom[140][101] = 16'h0048;
        rom[140][102] = 16'hFFF6;
        rom[140][103] = 16'h000F;
        rom[140][104] = 16'h000A;
        rom[140][105] = 16'h000A;
        rom[140][106] = 16'hFFF5;
        rom[140][107] = 16'hFFEB;
        rom[140][108] = 16'hFFF4;
        rom[140][109] = 16'h0026;
        rom[140][110] = 16'hFFD2;
        rom[140][111] = 16'hFFEF;
        rom[140][112] = 16'h0024;
        rom[140][113] = 16'hFFEC;
        rom[140][114] = 16'hFFFC;
        rom[140][115] = 16'hFFEA;
        rom[140][116] = 16'h0021;
        rom[140][117] = 16'h0021;
        rom[140][118] = 16'hFFDE;
        rom[140][119] = 16'hFFC8;
        rom[140][120] = 16'h0029;
        rom[140][121] = 16'h0011;
        rom[140][122] = 16'hFFF8;
        rom[140][123] = 16'h0038;
        rom[140][124] = 16'hFFF1;
        rom[140][125] = 16'hFFF7;
        rom[140][126] = 16'hFFE2;
        rom[140][127] = 16'h0027;
        rom[141][0] = 16'h0007;
        rom[141][1] = 16'hFFD0;
        rom[141][2] = 16'hFFFC;
        rom[141][3] = 16'h0016;
        rom[141][4] = 16'hFFDB;
        rom[141][5] = 16'h0018;
        rom[141][6] = 16'h0004;
        rom[141][7] = 16'hFFCA;
        rom[141][8] = 16'hFFF6;
        rom[141][9] = 16'hFFF6;
        rom[141][10] = 16'hFFEA;
        rom[141][11] = 16'h000C;
        rom[141][12] = 16'h001D;
        rom[141][13] = 16'hFFEF;
        rom[141][14] = 16'h0010;
        rom[141][15] = 16'hFFE4;
        rom[141][16] = 16'hFFF4;
        rom[141][17] = 16'hFFD5;
        rom[141][18] = 16'h0003;
        rom[141][19] = 16'h0008;
        rom[141][20] = 16'h0017;
        rom[141][21] = 16'hFFBD;
        rom[141][22] = 16'hFFF9;
        rom[141][23] = 16'h0006;
        rom[141][24] = 16'hFFEE;
        rom[141][25] = 16'h0028;
        rom[141][26] = 16'hFFDC;
        rom[141][27] = 16'h001B;
        rom[141][28] = 16'hFFEB;
        rom[141][29] = 16'hFFEC;
        rom[141][30] = 16'hFFEA;
        rom[141][31] = 16'hFFD4;
        rom[141][32] = 16'h0012;
        rom[141][33] = 16'hFFCE;
        rom[141][34] = 16'hFFF6;
        rom[141][35] = 16'h0021;
        rom[141][36] = 16'h000A;
        rom[141][37] = 16'h0011;
        rom[141][38] = 16'hFFE0;
        rom[141][39] = 16'hFFFD;
        rom[141][40] = 16'hFFAC;
        rom[141][41] = 16'hFFDB;
        rom[141][42] = 16'h0028;
        rom[141][43] = 16'hFFEE;
        rom[141][44] = 16'hFFE8;
        rom[141][45] = 16'h0013;
        rom[141][46] = 16'hFFE5;
        rom[141][47] = 16'h000F;
        rom[141][48] = 16'h0022;
        rom[141][49] = 16'h003A;
        rom[141][50] = 16'h002E;
        rom[141][51] = 16'h0017;
        rom[141][52] = 16'hFFF0;
        rom[141][53] = 16'hFFE4;
        rom[141][54] = 16'hFFE0;
        rom[141][55] = 16'hFFF5;
        rom[141][56] = 16'hFFF1;
        rom[141][57] = 16'hFFE4;
        rom[141][58] = 16'hFFD6;
        rom[141][59] = 16'h0024;
        rom[141][60] = 16'h0007;
        rom[141][61] = 16'h0013;
        rom[141][62] = 16'h0024;
        rom[141][63] = 16'hFFF7;
        rom[141][64] = 16'hFFF9;
        rom[141][65] = 16'hFFDB;
        rom[141][66] = 16'h0010;
        rom[141][67] = 16'h0009;
        rom[141][68] = 16'h0033;
        rom[141][69] = 16'h000C;
        rom[141][70] = 16'hFFE6;
        rom[141][71] = 16'hFFFB;
        rom[141][72] = 16'h0000;
        rom[141][73] = 16'hFFEC;
        rom[141][74] = 16'hFFC6;
        rom[141][75] = 16'hFFF3;
        rom[141][76] = 16'hFFFB;
        rom[141][77] = 16'hFFEA;
        rom[141][78] = 16'hFFF2;
        rom[141][79] = 16'hFFE3;
        rom[141][80] = 16'h003B;
        rom[141][81] = 16'h001B;
        rom[141][82] = 16'h0038;
        rom[141][83] = 16'hFFEB;
        rom[141][84] = 16'h0011;
        rom[141][85] = 16'hFFEF;
        rom[141][86] = 16'hFFDB;
        rom[141][87] = 16'hFFF1;
        rom[141][88] = 16'hFFEC;
        rom[141][89] = 16'h000B;
        rom[141][90] = 16'hFFFF;
        rom[141][91] = 16'h0016;
        rom[141][92] = 16'h0041;
        rom[141][93] = 16'h0014;
        rom[141][94] = 16'hFFE1;
        rom[141][95] = 16'h0038;
        rom[141][96] = 16'h0002;
        rom[141][97] = 16'h0017;
        rom[141][98] = 16'h000E;
        rom[141][99] = 16'hFFFB;
        rom[141][100] = 16'h0007;
        rom[141][101] = 16'hFFE1;
        rom[141][102] = 16'h0008;
        rom[141][103] = 16'h001B;
        rom[141][104] = 16'h000A;
        rom[141][105] = 16'hFFDE;
        rom[141][106] = 16'h0024;
        rom[141][107] = 16'h0027;
        rom[141][108] = 16'h002B;
        rom[141][109] = 16'h0024;
        rom[141][110] = 16'h0026;
        rom[141][111] = 16'h0016;
        rom[141][112] = 16'h0023;
        rom[141][113] = 16'hFFD7;
        rom[141][114] = 16'h0023;
        rom[141][115] = 16'hFFD7;
        rom[141][116] = 16'hFFD9;
        rom[141][117] = 16'h000E;
        rom[141][118] = 16'hFFE5;
        rom[141][119] = 16'h0008;
        rom[141][120] = 16'hFFFE;
        rom[141][121] = 16'h002A;
        rom[141][122] = 16'h0001;
        rom[141][123] = 16'h004B;
        rom[141][124] = 16'hFFEC;
        rom[141][125] = 16'hFFED;
        rom[141][126] = 16'h0002;
        rom[141][127] = 16'hFFF4;
        rom[142][0] = 16'h0025;
        rom[142][1] = 16'hFFD5;
        rom[142][2] = 16'h0013;
        rom[142][3] = 16'h0031;
        rom[142][4] = 16'hFFCF;
        rom[142][5] = 16'hFFED;
        rom[142][6] = 16'hFFE6;
        rom[142][7] = 16'hFFE5;
        rom[142][8] = 16'hFFDF;
        rom[142][9] = 16'h0028;
        rom[142][10] = 16'h0005;
        rom[142][11] = 16'h000A;
        rom[142][12] = 16'h0035;
        rom[142][13] = 16'hFFFE;
        rom[142][14] = 16'hFFD2;
        rom[142][15] = 16'h0012;
        rom[142][16] = 16'h0005;
        rom[142][17] = 16'hFFDE;
        rom[142][18] = 16'hFFFA;
        rom[142][19] = 16'hFFFB;
        rom[142][20] = 16'hFFF1;
        rom[142][21] = 16'h0008;
        rom[142][22] = 16'h000A;
        rom[142][23] = 16'hFFC3;
        rom[142][24] = 16'h0005;
        rom[142][25] = 16'hFFCE;
        rom[142][26] = 16'hFFFF;
        rom[142][27] = 16'hFFEE;
        rom[142][28] = 16'hFFE0;
        rom[142][29] = 16'h0014;
        rom[142][30] = 16'hFFEC;
        rom[142][31] = 16'h000D;
        rom[142][32] = 16'h000E;
        rom[142][33] = 16'hFFD3;
        rom[142][34] = 16'hFFF0;
        rom[142][35] = 16'h0002;
        rom[142][36] = 16'hFFE9;
        rom[142][37] = 16'hFFF7;
        rom[142][38] = 16'h002E;
        rom[142][39] = 16'h0001;
        rom[142][40] = 16'h0009;
        rom[142][41] = 16'hFFE5;
        rom[142][42] = 16'h0026;
        rom[142][43] = 16'hFFDE;
        rom[142][44] = 16'h003D;
        rom[142][45] = 16'h001E;
        rom[142][46] = 16'hFFFC;
        rom[142][47] = 16'hFFD8;
        rom[142][48] = 16'hFFFC;
        rom[142][49] = 16'hFFBB;
        rom[142][50] = 16'h0015;
        rom[142][51] = 16'h0004;
        rom[142][52] = 16'hFFF9;
        rom[142][53] = 16'h001A;
        rom[142][54] = 16'hFFF3;
        rom[142][55] = 16'h000B;
        rom[142][56] = 16'hFFFE;
        rom[142][57] = 16'hFFF4;
        rom[142][58] = 16'hFFDF;
        rom[142][59] = 16'h000A;
        rom[142][60] = 16'h0009;
        rom[142][61] = 16'h001E;
        rom[142][62] = 16'hFFCE;
        rom[142][63] = 16'hFFB6;
        rom[142][64] = 16'hFFF9;
        rom[142][65] = 16'h001E;
        rom[142][66] = 16'hFFD3;
        rom[142][67] = 16'h0002;
        rom[142][68] = 16'hFFC5;
        rom[142][69] = 16'hFFE7;
        rom[142][70] = 16'hFFFD;
        rom[142][71] = 16'hFFFB;
        rom[142][72] = 16'h002A;
        rom[142][73] = 16'h0003;
        rom[142][74] = 16'hFFF2;
        rom[142][75] = 16'hFFF9;
        rom[142][76] = 16'h0002;
        rom[142][77] = 16'hFFEB;
        rom[142][78] = 16'hFFE5;
        rom[142][79] = 16'h002F;
        rom[142][80] = 16'hFFD9;
        rom[142][81] = 16'hFFE5;
        rom[142][82] = 16'hFFC6;
        rom[142][83] = 16'h0024;
        rom[142][84] = 16'h0023;
        rom[142][85] = 16'h0011;
        rom[142][86] = 16'h0028;
        rom[142][87] = 16'h001B;
        rom[142][88] = 16'h0007;
        rom[142][89] = 16'h000B;
        rom[142][90] = 16'h0010;
        rom[142][91] = 16'h0021;
        rom[142][92] = 16'hFFFA;
        rom[142][93] = 16'hFFDA;
        rom[142][94] = 16'h0012;
        rom[142][95] = 16'h0017;
        rom[142][96] = 16'hFFCB;
        rom[142][97] = 16'hFFC5;
        rom[142][98] = 16'hFFDC;
        rom[142][99] = 16'hFFEB;
        rom[142][100] = 16'hFFFC;
        rom[142][101] = 16'h0013;
        rom[142][102] = 16'hFFC7;
        rom[142][103] = 16'hFFB9;
        rom[142][104] = 16'h000C;
        rom[142][105] = 16'hFFD2;
        rom[142][106] = 16'hFFE5;
        rom[142][107] = 16'h0002;
        rom[142][108] = 16'h0021;
        rom[142][109] = 16'hFFCF;
        rom[142][110] = 16'h0001;
        rom[142][111] = 16'hFFF4;
        rom[142][112] = 16'hFFDC;
        rom[142][113] = 16'hFFE9;
        rom[142][114] = 16'hFFD4;
        rom[142][115] = 16'h001D;
        rom[142][116] = 16'hFFE1;
        rom[142][117] = 16'hFFCE;
        rom[142][118] = 16'hFFC5;
        rom[142][119] = 16'hFFF8;
        rom[142][120] = 16'h0029;
        rom[142][121] = 16'hFFE1;
        rom[142][122] = 16'hFFFD;
        rom[142][123] = 16'h0002;
        rom[142][124] = 16'h0024;
        rom[142][125] = 16'h0003;
        rom[142][126] = 16'h0007;
        rom[142][127] = 16'h0019;
        rom[143][0] = 16'h0023;
        rom[143][1] = 16'h0000;
        rom[143][2] = 16'hFFD0;
        rom[143][3] = 16'h0015;
        rom[143][4] = 16'h000B;
        rom[143][5] = 16'hFFE5;
        rom[143][6] = 16'hFFDD;
        rom[143][7] = 16'hFFF8;
        rom[143][8] = 16'hFFF2;
        rom[143][9] = 16'hFFF0;
        rom[143][10] = 16'hFFF5;
        rom[143][11] = 16'hFFC3;
        rom[143][12] = 16'h0000;
        rom[143][13] = 16'h000C;
        rom[143][14] = 16'hFFEE;
        rom[143][15] = 16'hFFDB;
        rom[143][16] = 16'hFFF6;
        rom[143][17] = 16'hFFF9;
        rom[143][18] = 16'h000A;
        rom[143][19] = 16'hFFD7;
        rom[143][20] = 16'h000C;
        rom[143][21] = 16'hFFEC;
        rom[143][22] = 16'hFFFD;
        rom[143][23] = 16'hFFCA;
        rom[143][24] = 16'hFFE3;
        rom[143][25] = 16'h0009;
        rom[143][26] = 16'h0013;
        rom[143][27] = 16'h0014;
        rom[143][28] = 16'h0007;
        rom[143][29] = 16'h000E;
        rom[143][30] = 16'h000B;
        rom[143][31] = 16'h000C;
        rom[143][32] = 16'hFFE1;
        rom[143][33] = 16'hFFB0;
        rom[143][34] = 16'hFFED;
        rom[143][35] = 16'hFFFE;
        rom[143][36] = 16'hFFE3;
        rom[143][37] = 16'hFFFE;
        rom[143][38] = 16'hFFBB;
        rom[143][39] = 16'hFFD9;
        rom[143][40] = 16'h0004;
        rom[143][41] = 16'h001E;
        rom[143][42] = 16'hFFF4;
        rom[143][43] = 16'hFFDB;
        rom[143][44] = 16'h000E;
        rom[143][45] = 16'h0024;
        rom[143][46] = 16'hFFE4;
        rom[143][47] = 16'h001C;
        rom[143][48] = 16'hFFC8;
        rom[143][49] = 16'hFFF2;
        rom[143][50] = 16'hFFD7;
        rom[143][51] = 16'h001F;
        rom[143][52] = 16'h001F;
        rom[143][53] = 16'h001B;
        rom[143][54] = 16'h0016;
        rom[143][55] = 16'hFFFB;
        rom[143][56] = 16'h0012;
        rom[143][57] = 16'hFFB7;
        rom[143][58] = 16'hFFE1;
        rom[143][59] = 16'h000B;
        rom[143][60] = 16'hFFFD;
        rom[143][61] = 16'hFFFD;
        rom[143][62] = 16'h0021;
        rom[143][63] = 16'hFFE1;
        rom[143][64] = 16'h0011;
        rom[143][65] = 16'h002C;
        rom[143][66] = 16'h000F;
        rom[143][67] = 16'hFFF9;
        rom[143][68] = 16'h001F;
        rom[143][69] = 16'h000E;
        rom[143][70] = 16'hFFCC;
        rom[143][71] = 16'h002D;
        rom[143][72] = 16'hFFED;
        rom[143][73] = 16'h0002;
        rom[143][74] = 16'h0004;
        rom[143][75] = 16'hFFC2;
        rom[143][76] = 16'h0064;
        rom[143][77] = 16'hFFEB;
        rom[143][78] = 16'h000E;
        rom[143][79] = 16'hFFE7;
        rom[143][80] = 16'h0016;
        rom[143][81] = 16'h000F;
        rom[143][82] = 16'hFFCC;
        rom[143][83] = 16'hFFFE;
        rom[143][84] = 16'hFFE9;
        rom[143][85] = 16'hFFDB;
        rom[143][86] = 16'hFFE1;
        rom[143][87] = 16'h0002;
        rom[143][88] = 16'h001E;
        rom[143][89] = 16'h000C;
        rom[143][90] = 16'hFFE8;
        rom[143][91] = 16'h001C;
        rom[143][92] = 16'h0013;
        rom[143][93] = 16'hFFFE;
        rom[143][94] = 16'h0002;
        rom[143][95] = 16'h0007;
        rom[143][96] = 16'h001E;
        rom[143][97] = 16'hFFF2;
        rom[143][98] = 16'h0002;
        rom[143][99] = 16'h0008;
        rom[143][100] = 16'hFFF0;
        rom[143][101] = 16'hFFDB;
        rom[143][102] = 16'hFFF4;
        rom[143][103] = 16'h0007;
        rom[143][104] = 16'h001B;
        rom[143][105] = 16'hFFF4;
        rom[143][106] = 16'hFFF1;
        rom[143][107] = 16'h0019;
        rom[143][108] = 16'hFFFE;
        rom[143][109] = 16'h0028;
        rom[143][110] = 16'hFFC5;
        rom[143][111] = 16'hFFF6;
        rom[143][112] = 16'hFFE9;
        rom[143][113] = 16'hFFD9;
        rom[143][114] = 16'h001B;
        rom[143][115] = 16'h001B;
        rom[143][116] = 16'hFFC1;
        rom[143][117] = 16'h0003;
        rom[143][118] = 16'h000C;
        rom[143][119] = 16'h0015;
        rom[143][120] = 16'h0017;
        rom[143][121] = 16'hFFF8;
        rom[143][122] = 16'h0000;
        rom[143][123] = 16'h0040;
        rom[143][124] = 16'h0004;
        rom[143][125] = 16'hFFFA;
        rom[143][126] = 16'h001F;
        rom[143][127] = 16'h0003;
        rom[144][0] = 16'hFFEA;
        rom[144][1] = 16'h0029;
        rom[144][2] = 16'h0003;
        rom[144][3] = 16'hFFE3;
        rom[144][4] = 16'h0027;
        rom[144][5] = 16'hFFBB;
        rom[144][6] = 16'h0001;
        rom[144][7] = 16'h0006;
        rom[144][8] = 16'hFFCD;
        rom[144][9] = 16'hFFFA;
        rom[144][10] = 16'hFFCD;
        rom[144][11] = 16'h0009;
        rom[144][12] = 16'h0012;
        rom[144][13] = 16'h001F;
        rom[144][14] = 16'hFFC0;
        rom[144][15] = 16'hFFE1;
        rom[144][16] = 16'hFFF0;
        rom[144][17] = 16'hFFF2;
        rom[144][18] = 16'hFFD5;
        rom[144][19] = 16'hFFE9;
        rom[144][20] = 16'h000D;
        rom[144][21] = 16'h000C;
        rom[144][22] = 16'hFFDD;
        rom[144][23] = 16'hFFEF;
        rom[144][24] = 16'h000F;
        rom[144][25] = 16'hFFBC;
        rom[144][26] = 16'h001B;
        rom[144][27] = 16'hFFE1;
        rom[144][28] = 16'hFFF7;
        rom[144][29] = 16'h0015;
        rom[144][30] = 16'h0009;
        rom[144][31] = 16'h000E;
        rom[144][32] = 16'hFFC7;
        rom[144][33] = 16'hFFD7;
        rom[144][34] = 16'h0017;
        rom[144][35] = 16'h0015;
        rom[144][36] = 16'h0011;
        rom[144][37] = 16'hFFF5;
        rom[144][38] = 16'hFFDC;
        rom[144][39] = 16'h000C;
        rom[144][40] = 16'h001D;
        rom[144][41] = 16'h0007;
        rom[144][42] = 16'h0012;
        rom[144][43] = 16'hFFF8;
        rom[144][44] = 16'h000D;
        rom[144][45] = 16'h0000;
        rom[144][46] = 16'h0015;
        rom[144][47] = 16'hFFF1;
        rom[144][48] = 16'hFFDE;
        rom[144][49] = 16'hFFFA;
        rom[144][50] = 16'hFFE5;
        rom[144][51] = 16'hFFDC;
        rom[144][52] = 16'hFFD9;
        rom[144][53] = 16'hFFF9;
        rom[144][54] = 16'h0027;
        rom[144][55] = 16'hFFE7;
        rom[144][56] = 16'hFFEA;
        rom[144][57] = 16'hFFE7;
        rom[144][58] = 16'h000E;
        rom[144][59] = 16'h0010;
        rom[144][60] = 16'h0002;
        rom[144][61] = 16'hFFF5;
        rom[144][62] = 16'h001B;
        rom[144][63] = 16'hFFB9;
        rom[144][64] = 16'hFFFC;
        rom[144][65] = 16'h0028;
        rom[144][66] = 16'hFFFF;
        rom[144][67] = 16'h0007;
        rom[144][68] = 16'h0022;
        rom[144][69] = 16'h003F;
        rom[144][70] = 16'hFFE1;
        rom[144][71] = 16'hFFFA;
        rom[144][72] = 16'hFFF4;
        rom[144][73] = 16'h0019;
        rom[144][74] = 16'h0033;
        rom[144][75] = 16'hFFE9;
        rom[144][76] = 16'h000D;
        rom[144][77] = 16'hFFFF;
        rom[144][78] = 16'h0024;
        rom[144][79] = 16'h0021;
        rom[144][80] = 16'h0028;
        rom[144][81] = 16'h0012;
        rom[144][82] = 16'hFFE1;
        rom[144][83] = 16'h0004;
        rom[144][84] = 16'h0011;
        rom[144][85] = 16'hFFF7;
        rom[144][86] = 16'hFFF4;
        rom[144][87] = 16'hFFFA;
        rom[144][88] = 16'h0012;
        rom[144][89] = 16'hFFE1;
        rom[144][90] = 16'hFFD2;
        rom[144][91] = 16'hFFF5;
        rom[144][92] = 16'hFFFC;
        rom[144][93] = 16'h000C;
        rom[144][94] = 16'h002C;
        rom[144][95] = 16'hFFEF;
        rom[144][96] = 16'h001C;
        rom[144][97] = 16'h000F;
        rom[144][98] = 16'h0035;
        rom[144][99] = 16'h0016;
        rom[144][100] = 16'hFFFC;
        rom[144][101] = 16'h0002;
        rom[144][102] = 16'hFFF3;
        rom[144][103] = 16'h000F;
        rom[144][104] = 16'hFFE2;
        rom[144][105] = 16'hFFBA;
        rom[144][106] = 16'hFFE0;
        rom[144][107] = 16'h0009;
        rom[144][108] = 16'hFFFD;
        rom[144][109] = 16'hFFFE;
        rom[144][110] = 16'hFFF5;
        rom[144][111] = 16'h0022;
        rom[144][112] = 16'h001E;
        rom[144][113] = 16'hFFCB;
        rom[144][114] = 16'h0001;
        rom[144][115] = 16'h0008;
        rom[144][116] = 16'h0007;
        rom[144][117] = 16'hFFD3;
        rom[144][118] = 16'hFFC9;
        rom[144][119] = 16'h0011;
        rom[144][120] = 16'hFFF4;
        rom[144][121] = 16'hFFD8;
        rom[144][122] = 16'h0007;
        rom[144][123] = 16'hFFB5;
        rom[144][124] = 16'h0012;
        rom[144][125] = 16'hFFE7;
        rom[144][126] = 16'hFFE3;
        rom[144][127] = 16'hFFD2;
        rom[145][0] = 16'hFFD0;
        rom[145][1] = 16'hFFF3;
        rom[145][2] = 16'hFFEF;
        rom[145][3] = 16'hFFFC;
        rom[145][4] = 16'hFFEA;
        rom[145][5] = 16'hFFCD;
        rom[145][6] = 16'h000F;
        rom[145][7] = 16'h0010;
        rom[145][8] = 16'h000B;
        rom[145][9] = 16'hFFB3;
        rom[145][10] = 16'hFFD8;
        rom[145][11] = 16'hFFF6;
        rom[145][12] = 16'hFFE1;
        rom[145][13] = 16'h000A;
        rom[145][14] = 16'h0007;
        rom[145][15] = 16'h0026;
        rom[145][16] = 16'h0011;
        rom[145][17] = 16'hFFD8;
        rom[145][18] = 16'h0019;
        rom[145][19] = 16'h0010;
        rom[145][20] = 16'hFFC8;
        rom[145][21] = 16'h0010;
        rom[145][22] = 16'h0004;
        rom[145][23] = 16'hFFF5;
        rom[145][24] = 16'hFFF3;
        rom[145][25] = 16'hFFFC;
        rom[145][26] = 16'hFFFE;
        rom[145][27] = 16'h0012;
        rom[145][28] = 16'h0021;
        rom[145][29] = 16'h0000;
        rom[145][30] = 16'hFFDF;
        rom[145][31] = 16'h000F;
        rom[145][32] = 16'hFFB1;
        rom[145][33] = 16'hFFF4;
        rom[145][34] = 16'h002E;
        rom[145][35] = 16'h0016;
        rom[145][36] = 16'h0023;
        rom[145][37] = 16'hFFE0;
        rom[145][38] = 16'hFFB5;
        rom[145][39] = 16'h0016;
        rom[145][40] = 16'hFFF8;
        rom[145][41] = 16'h001A;
        rom[145][42] = 16'hFFCB;
        rom[145][43] = 16'hFFFE;
        rom[145][44] = 16'hFFF0;
        rom[145][45] = 16'h0032;
        rom[145][46] = 16'h0011;
        rom[145][47] = 16'hFFD6;
        rom[145][48] = 16'h0002;
        rom[145][49] = 16'h0005;
        rom[145][50] = 16'hFFD9;
        rom[145][51] = 16'hFFBD;
        rom[145][52] = 16'h0041;
        rom[145][53] = 16'hFFFD;
        rom[145][54] = 16'hFFF9;
        rom[145][55] = 16'h001E;
        rom[145][56] = 16'h0000;
        rom[145][57] = 16'hFFE7;
        rom[145][58] = 16'hFFD0;
        rom[145][59] = 16'hFFCD;
        rom[145][60] = 16'hFFF5;
        rom[145][61] = 16'h0008;
        rom[145][62] = 16'h001A;
        rom[145][63] = 16'h0007;
        rom[145][64] = 16'h0009;
        rom[145][65] = 16'h0007;
        rom[145][66] = 16'hFFE9;
        rom[145][67] = 16'hFFF0;
        rom[145][68] = 16'h0009;
        rom[145][69] = 16'h001B;
        rom[145][70] = 16'hFFD3;
        rom[145][71] = 16'hFFFA;
        rom[145][72] = 16'hFFD5;
        rom[145][73] = 16'hFFDF;
        rom[145][74] = 16'hFFEF;
        rom[145][75] = 16'hFFE1;
        rom[145][76] = 16'hFFF0;
        rom[145][77] = 16'hFFBA;
        rom[145][78] = 16'h0008;
        rom[145][79] = 16'hFFE1;
        rom[145][80] = 16'h000D;
        rom[145][81] = 16'h001F;
        rom[145][82] = 16'hFFDD;
        rom[145][83] = 16'hFFEF;
        rom[145][84] = 16'h0010;
        rom[145][85] = 16'hFFED;
        rom[145][86] = 16'h001D;
        rom[145][87] = 16'hFFD9;
        rom[145][88] = 16'hFFE8;
        rom[145][89] = 16'h0002;
        rom[145][90] = 16'hFFCA;
        rom[145][91] = 16'h0005;
        rom[145][92] = 16'hFFE6;
        rom[145][93] = 16'h0008;
        rom[145][94] = 16'hFFDF;
        rom[145][95] = 16'hFFF9;
        rom[145][96] = 16'hFFE4;
        rom[145][97] = 16'hFFEF;
        rom[145][98] = 16'h0014;
        rom[145][99] = 16'hFFEF;
        rom[145][100] = 16'h002F;
        rom[145][101] = 16'hFFFA;
        rom[145][102] = 16'h0000;
        rom[145][103] = 16'h0002;
        rom[145][104] = 16'hFFBE;
        rom[145][105] = 16'hFFD3;
        rom[145][106] = 16'hFFED;
        rom[145][107] = 16'h000A;
        rom[145][108] = 16'hFFEA;
        rom[145][109] = 16'h000C;
        rom[145][110] = 16'hFFD7;
        rom[145][111] = 16'h000E;
        rom[145][112] = 16'hFFE8;
        rom[145][113] = 16'h001C;
        rom[145][114] = 16'h001F;
        rom[145][115] = 16'h0030;
        rom[145][116] = 16'h000C;
        rom[145][117] = 16'h0001;
        rom[145][118] = 16'hFFE2;
        rom[145][119] = 16'h0027;
        rom[145][120] = 16'hFFE1;
        rom[145][121] = 16'hFFF4;
        rom[145][122] = 16'h0002;
        rom[145][123] = 16'h000C;
        rom[145][124] = 16'h0008;
        rom[145][125] = 16'hFFB1;
        rom[145][126] = 16'h0008;
        rom[145][127] = 16'h001D;
        rom[146][0] = 16'h0014;
        rom[146][1] = 16'h000A;
        rom[146][2] = 16'h0036;
        rom[146][3] = 16'hFFE7;
        rom[146][4] = 16'h000A;
        rom[146][5] = 16'h000D;
        rom[146][6] = 16'h0025;
        rom[146][7] = 16'hFFC8;
        rom[146][8] = 16'hFFF6;
        rom[146][9] = 16'h0024;
        rom[146][10] = 16'h0007;
        rom[146][11] = 16'h0002;
        rom[146][12] = 16'hFFE0;
        rom[146][13] = 16'h0011;
        rom[146][14] = 16'hFFF0;
        rom[146][15] = 16'h0027;
        rom[146][16] = 16'h000D;
        rom[146][17] = 16'hFFCD;
        rom[146][18] = 16'hFFF3;
        rom[146][19] = 16'hFFFE;
        rom[146][20] = 16'hFFF9;
        rom[146][21] = 16'h0019;
        rom[146][22] = 16'h002B;
        rom[146][23] = 16'h0007;
        rom[146][24] = 16'h000C;
        rom[146][25] = 16'h001B;
        rom[146][26] = 16'hFFCF;
        rom[146][27] = 16'h0023;
        rom[146][28] = 16'h001A;
        rom[146][29] = 16'h000E;
        rom[146][30] = 16'h0004;
        rom[146][31] = 16'hFFA1;
        rom[146][32] = 16'hFFCD;
        rom[146][33] = 16'h0011;
        rom[146][34] = 16'hFFCB;
        rom[146][35] = 16'hFFF3;
        rom[146][36] = 16'hFFB6;
        rom[146][37] = 16'h0002;
        rom[146][38] = 16'h001E;
        rom[146][39] = 16'h001F;
        rom[146][40] = 16'hFFE6;
        rom[146][41] = 16'h0016;
        rom[146][42] = 16'hFFF1;
        rom[146][43] = 16'hFFF6;
        rom[146][44] = 16'hFFB9;
        rom[146][45] = 16'h0009;
        rom[146][46] = 16'h0009;
        rom[146][47] = 16'h0008;
        rom[146][48] = 16'hFFE4;
        rom[146][49] = 16'h0015;
        rom[146][50] = 16'h0017;
        rom[146][51] = 16'h0015;
        rom[146][52] = 16'h001B;
        rom[146][53] = 16'hFFB2;
        rom[146][54] = 16'hFFE3;
        rom[146][55] = 16'hFFEC;
        rom[146][56] = 16'hFFD0;
        rom[146][57] = 16'hFFCA;
        rom[146][58] = 16'hFFB6;
        rom[146][59] = 16'hFFDF;
        rom[146][60] = 16'hFFEF;
        rom[146][61] = 16'h0007;
        rom[146][62] = 16'h001C;
        rom[146][63] = 16'hFFD7;
        rom[146][64] = 16'h0013;
        rom[146][65] = 16'hFFDE;
        rom[146][66] = 16'hFFF8;
        rom[146][67] = 16'hFFF9;
        rom[146][68] = 16'h000C;
        rom[146][69] = 16'hFFF9;
        rom[146][70] = 16'h0016;
        rom[146][71] = 16'h000A;
        rom[146][72] = 16'hFFE5;
        rom[146][73] = 16'h0035;
        rom[146][74] = 16'hFFDF;
        rom[146][75] = 16'h000A;
        rom[146][76] = 16'h000C;
        rom[146][77] = 16'hFFFE;
        rom[146][78] = 16'hFFEF;
        rom[146][79] = 16'hFFFB;
        rom[146][80] = 16'h000E;
        rom[146][81] = 16'hFFFD;
        rom[146][82] = 16'h000A;
        rom[146][83] = 16'hFFDC;
        rom[146][84] = 16'hFFC8;
        rom[146][85] = 16'hFFEE;
        rom[146][86] = 16'h000D;
        rom[146][87] = 16'hFFFA;
        rom[146][88] = 16'hFFC7;
        rom[146][89] = 16'hFFE9;
        rom[146][90] = 16'hFFEE;
        rom[146][91] = 16'hFFF0;
        rom[146][92] = 16'h000C;
        rom[146][93] = 16'hFFF6;
        rom[146][94] = 16'hFFCE;
        rom[146][95] = 16'h0015;
        rom[146][96] = 16'hFFFE;
        rom[146][97] = 16'hFFFD;
        rom[146][98] = 16'h000F;
        rom[146][99] = 16'hFFEF;
        rom[146][100] = 16'h0009;
        rom[146][101] = 16'h001A;
        rom[146][102] = 16'h002F;
        rom[146][103] = 16'h0025;
        rom[146][104] = 16'hFFFB;
        rom[146][105] = 16'hFFCC;
        rom[146][106] = 16'hFFF1;
        rom[146][107] = 16'hFFEC;
        rom[146][108] = 16'h001D;
        rom[146][109] = 16'h0033;
        rom[146][110] = 16'h0012;
        rom[146][111] = 16'hFFFE;
        rom[146][112] = 16'h0016;
        rom[146][113] = 16'h0005;
        rom[146][114] = 16'h001F;
        rom[146][115] = 16'hFFE1;
        rom[146][116] = 16'h0029;
        rom[146][117] = 16'h000A;
        rom[146][118] = 16'h0008;
        rom[146][119] = 16'hFFF9;
        rom[146][120] = 16'h0011;
        rom[146][121] = 16'h000B;
        rom[146][122] = 16'h001C;
        rom[146][123] = 16'h0006;
        rom[146][124] = 16'hFFDB;
        rom[146][125] = 16'h000C;
        rom[146][126] = 16'h0016;
        rom[146][127] = 16'hFFE4;
        rom[147][0] = 16'hFFC8;
        rom[147][1] = 16'h0012;
        rom[147][2] = 16'h0000;
        rom[147][3] = 16'hFFD3;
        rom[147][4] = 16'h0026;
        rom[147][5] = 16'h0033;
        rom[147][6] = 16'h0030;
        rom[147][7] = 16'hFFD2;
        rom[147][8] = 16'hFFE8;
        rom[147][9] = 16'h001D;
        rom[147][10] = 16'hFFE2;
        rom[147][11] = 16'h001D;
        rom[147][12] = 16'h0019;
        rom[147][13] = 16'h0010;
        rom[147][14] = 16'h003E;
        rom[147][15] = 16'h0024;
        rom[147][16] = 16'hFFFE;
        rom[147][17] = 16'h000E;
        rom[147][18] = 16'hFFDC;
        rom[147][19] = 16'h0003;
        rom[147][20] = 16'h0009;
        rom[147][21] = 16'hFFE0;
        rom[147][22] = 16'hFFCB;
        rom[147][23] = 16'h001E;
        rom[147][24] = 16'hFFDC;
        rom[147][25] = 16'h0007;
        rom[147][26] = 16'h0011;
        rom[147][27] = 16'h001D;
        rom[147][28] = 16'hFFF1;
        rom[147][29] = 16'h000E;
        rom[147][30] = 16'hFFDF;
        rom[147][31] = 16'hFFE1;
        rom[147][32] = 16'h0001;
        rom[147][33] = 16'hFFD1;
        rom[147][34] = 16'h0009;
        rom[147][35] = 16'h0010;
        rom[147][36] = 16'hFFE9;
        rom[147][37] = 16'hFFF5;
        rom[147][38] = 16'h0011;
        rom[147][39] = 16'h0000;
        rom[147][40] = 16'hFFE2;
        rom[147][41] = 16'hFFFA;
        rom[147][42] = 16'hFFDC;
        rom[147][43] = 16'hFFAB;
        rom[147][44] = 16'hFFEE;
        rom[147][45] = 16'hFFE1;
        rom[147][46] = 16'h0004;
        rom[147][47] = 16'hFFFA;
        rom[147][48] = 16'h0010;
        rom[147][49] = 16'hFFFE;
        rom[147][50] = 16'h0042;
        rom[147][51] = 16'hFFEB;
        rom[147][52] = 16'hFFF3;
        rom[147][53] = 16'hFFD8;
        rom[147][54] = 16'h0023;
        rom[147][55] = 16'hFFF9;
        rom[147][56] = 16'h0006;
        rom[147][57] = 16'hFFD7;
        rom[147][58] = 16'hFFE6;
        rom[147][59] = 16'h001D;
        rom[147][60] = 16'hFFFA;
        rom[147][61] = 16'h0028;
        rom[147][62] = 16'h0000;
        rom[147][63] = 16'h0015;
        rom[147][64] = 16'hFFDD;
        rom[147][65] = 16'hFFC9;
        rom[147][66] = 16'h001A;
        rom[147][67] = 16'h0035;
        rom[147][68] = 16'h000C;
        rom[147][69] = 16'h0029;
        rom[147][70] = 16'h001B;
        rom[147][71] = 16'hFFC8;
        rom[147][72] = 16'hFFE9;
        rom[147][73] = 16'h0027;
        rom[147][74] = 16'hFFD1;
        rom[147][75] = 16'h0003;
        rom[147][76] = 16'h0009;
        rom[147][77] = 16'hFFDF;
        rom[147][78] = 16'hFFF8;
        rom[147][79] = 16'hFFEB;
        rom[147][80] = 16'h0014;
        rom[147][81] = 16'h001E;
        rom[147][82] = 16'hFFFD;
        rom[147][83] = 16'hFFF4;
        rom[147][84] = 16'h000D;
        rom[147][85] = 16'h000B;
        rom[147][86] = 16'hFFE6;
        rom[147][87] = 16'hFFE7;
        rom[147][88] = 16'h0009;
        rom[147][89] = 16'h0005;
        rom[147][90] = 16'h0023;
        rom[147][91] = 16'hFFD2;
        rom[147][92] = 16'hFFF9;
        rom[147][93] = 16'h001B;
        rom[147][94] = 16'hFFD0;
        rom[147][95] = 16'hFFD5;
        rom[147][96] = 16'hFFF2;
        rom[147][97] = 16'h0002;
        rom[147][98] = 16'h002D;
        rom[147][99] = 16'hFFF2;
        rom[147][100] = 16'h0007;
        rom[147][101] = 16'hFFF8;
        rom[147][102] = 16'hFFF9;
        rom[147][103] = 16'hFFF2;
        rom[147][104] = 16'hFFCD;
        rom[147][105] = 16'hFFDC;
        rom[147][106] = 16'h0026;
        rom[147][107] = 16'h0023;
        rom[147][108] = 16'h0007;
        rom[147][109] = 16'h000E;
        rom[147][110] = 16'h002E;
        rom[147][111] = 16'h0014;
        rom[147][112] = 16'h001C;
        rom[147][113] = 16'hFFE4;
        rom[147][114] = 16'h0016;
        rom[147][115] = 16'hFFDF;
        rom[147][116] = 16'hFFE3;
        rom[147][117] = 16'h0020;
        rom[147][118] = 16'h0044;
        rom[147][119] = 16'h0028;
        rom[147][120] = 16'hFFD6;
        rom[147][121] = 16'h000E;
        rom[147][122] = 16'hFFF8;
        rom[147][123] = 16'hFFE5;
        rom[147][124] = 16'hFFF4;
        rom[147][125] = 16'hFFFE;
        rom[147][126] = 16'hFFE7;
        rom[147][127] = 16'hFFB9;
        rom[148][0] = 16'h0002;
        rom[148][1] = 16'hFFFD;
        rom[148][2] = 16'hFFC1;
        rom[148][3] = 16'h0025;
        rom[148][4] = 16'hFFE9;
        rom[148][5] = 16'hFFFE;
        rom[148][6] = 16'h0009;
        rom[148][7] = 16'hFFF2;
        rom[148][8] = 16'h001B;
        rom[148][9] = 16'h0016;
        rom[148][10] = 16'hFFBF;
        rom[148][11] = 16'hFFBE;
        rom[148][12] = 16'h000E;
        rom[148][13] = 16'hFFD5;
        rom[148][14] = 16'h000D;
        rom[148][15] = 16'hFFF4;
        rom[148][16] = 16'h0015;
        rom[148][17] = 16'hFFF3;
        rom[148][18] = 16'h0007;
        rom[148][19] = 16'hFFD2;
        rom[148][20] = 16'hFFBE;
        rom[148][21] = 16'h0003;
        rom[148][22] = 16'hFFAF;
        rom[148][23] = 16'hFFDC;
        rom[148][24] = 16'hFFFC;
        rom[148][25] = 16'hFFEF;
        rom[148][26] = 16'h0019;
        rom[148][27] = 16'hFFE7;
        rom[148][28] = 16'hFFDA;
        rom[148][29] = 16'hFFD1;
        rom[148][30] = 16'hFFEF;
        rom[148][31] = 16'h0001;
        rom[148][32] = 16'hFFBF;
        rom[148][33] = 16'hFFE7;
        rom[148][34] = 16'hFFEA;
        rom[148][35] = 16'hFFE5;
        rom[148][36] = 16'hFFFF;
        rom[148][37] = 16'hFFEA;
        rom[148][38] = 16'h000E;
        rom[148][39] = 16'h0018;
        rom[148][40] = 16'h000C;
        rom[148][41] = 16'h000C;
        rom[148][42] = 16'h001F;
        rom[148][43] = 16'h0016;
        rom[148][44] = 16'h000E;
        rom[148][45] = 16'hFFC9;
        rom[148][46] = 16'h000A;
        rom[148][47] = 16'h0012;
        rom[148][48] = 16'hFFF3;
        rom[148][49] = 16'h0005;
        rom[148][50] = 16'hFFF5;
        rom[148][51] = 16'h0008;
        rom[148][52] = 16'hFFF7;
        rom[148][53] = 16'hFFEC;
        rom[148][54] = 16'hFFF2;
        rom[148][55] = 16'hFFF5;
        rom[148][56] = 16'h000C;
        rom[148][57] = 16'h0010;
        rom[148][58] = 16'h0016;
        rom[148][59] = 16'hFFE5;
        rom[148][60] = 16'hFFFD;
        rom[148][61] = 16'hFFD7;
        rom[148][62] = 16'h0008;
        rom[148][63] = 16'hFFE3;
        rom[148][64] = 16'hFFFE;
        rom[148][65] = 16'h0001;
        rom[148][66] = 16'h000A;
        rom[148][67] = 16'h0015;
        rom[148][68] = 16'h000D;
        rom[148][69] = 16'hFFF4;
        rom[148][70] = 16'hFFEA;
        rom[148][71] = 16'hFFCA;
        rom[148][72] = 16'h0000;
        rom[148][73] = 16'h0006;
        rom[148][74] = 16'hFFEC;
        rom[148][75] = 16'hFFF9;
        rom[148][76] = 16'hFFD4;
        rom[148][77] = 16'h0017;
        rom[148][78] = 16'h0023;
        rom[148][79] = 16'h0013;
        rom[148][80] = 16'h0000;
        rom[148][81] = 16'hFFFF;
        rom[148][82] = 16'hFFE3;
        rom[148][83] = 16'hFFEA;
        rom[148][84] = 16'h000C;
        rom[148][85] = 16'hFFF7;
        rom[148][86] = 16'hFFD0;
        rom[148][87] = 16'h0004;
        rom[148][88] = 16'hFFC6;
        rom[148][89] = 16'h000C;
        rom[148][90] = 16'hFFEA;
        rom[148][91] = 16'h0030;
        rom[148][92] = 16'h0036;
        rom[148][93] = 16'hFFAB;
        rom[148][94] = 16'h0017;
        rom[148][95] = 16'hFFF6;
        rom[148][96] = 16'hFFF6;
        rom[148][97] = 16'h0016;
        rom[148][98] = 16'hFFDE;
        rom[148][99] = 16'hFFE2;
        rom[148][100] = 16'hFFC8;
        rom[148][101] = 16'h0007;
        rom[148][102] = 16'hFFCA;
        rom[148][103] = 16'hFFEB;
        rom[148][104] = 16'h000A;
        rom[148][105] = 16'hFFDC;
        rom[148][106] = 16'h002A;
        rom[148][107] = 16'hFFCF;
        rom[148][108] = 16'hFFC8;
        rom[148][109] = 16'hFFED;
        rom[148][110] = 16'hFFD5;
        rom[148][111] = 16'hFFF0;
        rom[148][112] = 16'hFFD2;
        rom[148][113] = 16'hFFEB;
        rom[148][114] = 16'hFFED;
        rom[148][115] = 16'h000C;
        rom[148][116] = 16'h0023;
        rom[148][117] = 16'h0021;
        rom[148][118] = 16'hFFF4;
        rom[148][119] = 16'hFFF8;
        rom[148][120] = 16'hFFE9;
        rom[148][121] = 16'hFFDA;
        rom[148][122] = 16'hFFF9;
        rom[148][123] = 16'h004B;
        rom[148][124] = 16'h000E;
        rom[148][125] = 16'h001E;
        rom[148][126] = 16'hFFE8;
        rom[148][127] = 16'hFFF0;
        rom[149][0] = 16'h0025;
        rom[149][1] = 16'h0006;
        rom[149][2] = 16'h0016;
        rom[149][3] = 16'h0007;
        rom[149][4] = 16'hFFE3;
        rom[149][5] = 16'hFFE4;
        rom[149][6] = 16'hFFC8;
        rom[149][7] = 16'h0025;
        rom[149][8] = 16'h0000;
        rom[149][9] = 16'h000B;
        rom[149][10] = 16'h0001;
        rom[149][11] = 16'hFFF6;
        rom[149][12] = 16'hFFF0;
        rom[149][13] = 16'hFFED;
        rom[149][14] = 16'h0018;
        rom[149][15] = 16'h000A;
        rom[149][16] = 16'hFFA2;
        rom[149][17] = 16'h002E;
        rom[149][18] = 16'h0007;
        rom[149][19] = 16'h0004;
        rom[149][20] = 16'h000F;
        rom[149][21] = 16'h0016;
        rom[149][22] = 16'hFFFA;
        rom[149][23] = 16'h0007;
        rom[149][24] = 16'h0011;
        rom[149][25] = 16'hFFC9;
        rom[149][26] = 16'h0019;
        rom[149][27] = 16'hFFE5;
        rom[149][28] = 16'hFFE5;
        rom[149][29] = 16'h0019;
        rom[149][30] = 16'hFFD7;
        rom[149][31] = 16'h0016;
        rom[149][32] = 16'h000C;
        rom[149][33] = 16'h000A;
        rom[149][34] = 16'hFFD2;
        rom[149][35] = 16'h0014;
        rom[149][36] = 16'hFFF5;
        rom[149][37] = 16'h0011;
        rom[149][38] = 16'h002C;
        rom[149][39] = 16'h001A;
        rom[149][40] = 16'hFFFD;
        rom[149][41] = 16'hFFFE;
        rom[149][42] = 16'hFFF6;
        rom[149][43] = 16'hFFDC;
        rom[149][44] = 16'hFFFB;
        rom[149][45] = 16'hFFFB;
        rom[149][46] = 16'h0004;
        rom[149][47] = 16'hFFDF;
        rom[149][48] = 16'h000D;
        rom[149][49] = 16'h0004;
        rom[149][50] = 16'h0016;
        rom[149][51] = 16'hFFE3;
        rom[149][52] = 16'hFFBB;
        rom[149][53] = 16'h0011;
        rom[149][54] = 16'hFFF9;
        rom[149][55] = 16'hFFC7;
        rom[149][56] = 16'h0007;
        rom[149][57] = 16'h0011;
        rom[149][58] = 16'hFFFB;
        rom[149][59] = 16'hFFFF;
        rom[149][60] = 16'hFFD5;
        rom[149][61] = 16'hFFFD;
        rom[149][62] = 16'hFFE1;
        rom[149][63] = 16'hFFE7;
        rom[149][64] = 16'h000A;
        rom[149][65] = 16'hFFF9;
        rom[149][66] = 16'h0005;
        rom[149][67] = 16'hFFEF;
        rom[149][68] = 16'hFFBD;
        rom[149][69] = 16'hFFD7;
        rom[149][70] = 16'h001D;
        rom[149][71] = 16'h0001;
        rom[149][72] = 16'hFFF8;
        rom[149][73] = 16'h0004;
        rom[149][74] = 16'hFFFD;
        rom[149][75] = 16'h0011;
        rom[149][76] = 16'hFFF6;
        rom[149][77] = 16'hFFD0;
        rom[149][78] = 16'h0003;
        rom[149][79] = 16'hFFC8;
        rom[149][80] = 16'h0006;
        rom[149][81] = 16'h0000;
        rom[149][82] = 16'h0009;
        rom[149][83] = 16'h0002;
        rom[149][84] = 16'h0015;
        rom[149][85] = 16'hFFD7;
        rom[149][86] = 16'h001D;
        rom[149][87] = 16'hFFD1;
        rom[149][88] = 16'h000A;
        rom[149][89] = 16'hFFCF;
        rom[149][90] = 16'h0007;
        rom[149][91] = 16'hFFDF;
        rom[149][92] = 16'h0003;
        rom[149][93] = 16'hFFAD;
        rom[149][94] = 16'hFFEE;
        rom[149][95] = 16'hFFE7;
        rom[149][96] = 16'hFF9B;
        rom[149][97] = 16'hFFCD;
        rom[149][98] = 16'hFFD8;
        rom[149][99] = 16'hFFDE;
        rom[149][100] = 16'hFFEA;
        rom[149][101] = 16'hFFF6;
        rom[149][102] = 16'hFFDE;
        rom[149][103] = 16'hFFFC;
        rom[149][104] = 16'hFFA4;
        rom[149][105] = 16'hFFB5;
        rom[149][106] = 16'h0007;
        rom[149][107] = 16'hFFF8;
        rom[149][108] = 16'h0012;
        rom[149][109] = 16'hFFD7;
        rom[149][110] = 16'hFFFE;
        rom[149][111] = 16'hFFC3;
        rom[149][112] = 16'hFFEA;
        rom[149][113] = 16'h0004;
        rom[149][114] = 16'hFFF4;
        rom[149][115] = 16'hFFF6;
        rom[149][116] = 16'hFFF4;
        rom[149][117] = 16'h0007;
        rom[149][118] = 16'hFFE9;
        rom[149][119] = 16'h000B;
        rom[149][120] = 16'hFFE1;
        rom[149][121] = 16'h000F;
        rom[149][122] = 16'hFFF9;
        rom[149][123] = 16'hFFD7;
        rom[149][124] = 16'hFFD1;
        rom[149][125] = 16'hFFD9;
        rom[149][126] = 16'hFFF3;
        rom[149][127] = 16'h000A;
        rom[150][0] = 16'hFFCF;
        rom[150][1] = 16'h0000;
        rom[150][2] = 16'hFFCA;
        rom[150][3] = 16'h000E;
        rom[150][4] = 16'h001F;
        rom[150][5] = 16'h0011;
        rom[150][6] = 16'hFFFE;
        rom[150][7] = 16'hFFFA;
        rom[150][8] = 16'h003D;
        rom[150][9] = 16'h0009;
        rom[150][10] = 16'hFFE6;
        rom[150][11] = 16'h0003;
        rom[150][12] = 16'h000B;
        rom[150][13] = 16'hFFFE;
        rom[150][14] = 16'h0006;
        rom[150][15] = 16'h001B;
        rom[150][16] = 16'h0019;
        rom[150][17] = 16'hFFF4;
        rom[150][18] = 16'h0009;
        rom[150][19] = 16'hFFE1;
        rom[150][20] = 16'hFFD0;
        rom[150][21] = 16'h0018;
        rom[150][22] = 16'hFFDC;
        rom[150][23] = 16'hFFDF;
        rom[150][24] = 16'hFFE5;
        rom[150][25] = 16'hFFF4;
        rom[150][26] = 16'h0029;
        rom[150][27] = 16'h0017;
        rom[150][28] = 16'hFFDC;
        rom[150][29] = 16'hFFB1;
        rom[150][30] = 16'h0022;
        rom[150][31] = 16'h0003;
        rom[150][32] = 16'hFFC2;
        rom[150][33] = 16'h000C;
        rom[150][34] = 16'hFFF5;
        rom[150][35] = 16'hFFD3;
        rom[150][36] = 16'h000E;
        rom[150][37] = 16'hFFEF;
        rom[150][38] = 16'hFFD3;
        rom[150][39] = 16'hFFFF;
        rom[150][40] = 16'h0016;
        rom[150][41] = 16'h0032;
        rom[150][42] = 16'h0007;
        rom[150][43] = 16'hFFF5;
        rom[150][44] = 16'h0005;
        rom[150][45] = 16'hFFCB;
        rom[150][46] = 16'hFFF4;
        rom[150][47] = 16'h000D;
        rom[150][48] = 16'hFFE5;
        rom[150][49] = 16'hFFDC;
        rom[150][50] = 16'hFFC8;
        rom[150][51] = 16'hFFEA;
        rom[150][52] = 16'hFFDB;
        rom[150][53] = 16'h0012;
        rom[150][54] = 16'h001B;
        rom[150][55] = 16'h0029;
        rom[150][56] = 16'hFFFD;
        rom[150][57] = 16'h000C;
        rom[150][58] = 16'h0010;
        rom[150][59] = 16'h0018;
        rom[150][60] = 16'h003A;
        rom[150][61] = 16'hFFDB;
        rom[150][62] = 16'hFFEF;
        rom[150][63] = 16'hFFE2;
        rom[150][64] = 16'hFFCD;
        rom[150][65] = 16'h001D;
        rom[150][66] = 16'hFFFC;
        rom[150][67] = 16'h001E;
        rom[150][68] = 16'h0000;
        rom[150][69] = 16'h0010;
        rom[150][70] = 16'h0015;
        rom[150][71] = 16'hFFB4;
        rom[150][72] = 16'hFFF1;
        rom[150][73] = 16'h0002;
        rom[150][74] = 16'hFFBE;
        rom[150][75] = 16'hFFEA;
        rom[150][76] = 16'hFFD1;
        rom[150][77] = 16'h001D;
        rom[150][78] = 16'h0027;
        rom[150][79] = 16'h0026;
        rom[150][80] = 16'hFFD9;
        rom[150][81] = 16'hFFFC;
        rom[150][82] = 16'hFFFB;
        rom[150][83] = 16'hFFF7;
        rom[150][84] = 16'h0011;
        rom[150][85] = 16'h0007;
        rom[150][86] = 16'hFFC3;
        rom[150][87] = 16'h000C;
        rom[150][88] = 16'hFFC8;
        rom[150][89] = 16'h0008;
        rom[150][90] = 16'hFFFB;
        rom[150][91] = 16'h0013;
        rom[150][92] = 16'hFFF9;
        rom[150][93] = 16'hFFAC;
        rom[150][94] = 16'hFFED;
        rom[150][95] = 16'h0000;
        rom[150][96] = 16'hFFEB;
        rom[150][97] = 16'h0000;
        rom[150][98] = 16'hFFDF;
        rom[150][99] = 16'hFFF4;
        rom[150][100] = 16'hFFC0;
        rom[150][101] = 16'hFFD4;
        rom[150][102] = 16'hFFC8;
        rom[150][103] = 16'hFFF3;
        rom[150][104] = 16'h0008;
        rom[150][105] = 16'hFFE0;
        rom[150][106] = 16'hFFF4;
        rom[150][107] = 16'hFFDC;
        rom[150][108] = 16'hFFE7;
        rom[150][109] = 16'hFFF4;
        rom[150][110] = 16'hFFFE;
        rom[150][111] = 16'h0006;
        rom[150][112] = 16'hFFC7;
        rom[150][113] = 16'h000D;
        rom[150][114] = 16'hFFEA;
        rom[150][115] = 16'h000D;
        rom[150][116] = 16'h000B;
        rom[150][117] = 16'h000F;
        rom[150][118] = 16'hFFF8;
        rom[150][119] = 16'hFFE0;
        rom[150][120] = 16'h000F;
        rom[150][121] = 16'hFFE9;
        rom[150][122] = 16'h0011;
        rom[150][123] = 16'h001A;
        rom[150][124] = 16'hFFFA;
        rom[150][125] = 16'h000E;
        rom[150][126] = 16'hFFD7;
        rom[150][127] = 16'h0000;
        rom[151][0] = 16'h002E;
        rom[151][1] = 16'hFFE5;
        rom[151][2] = 16'hFFDE;
        rom[151][3] = 16'h0006;
        rom[151][4] = 16'h0008;
        rom[151][5] = 16'hFFA4;
        rom[151][6] = 16'h0006;
        rom[151][7] = 16'h000C;
        rom[151][8] = 16'h0001;
        rom[151][9] = 16'hFFCF;
        rom[151][10] = 16'h001D;
        rom[151][11] = 16'hFFBF;
        rom[151][12] = 16'h0013;
        rom[151][13] = 16'hFFF4;
        rom[151][14] = 16'hFFEB;
        rom[151][15] = 16'h000C;
        rom[151][16] = 16'hFFD8;
        rom[151][17] = 16'hFFD0;
        rom[151][18] = 16'hFFF9;
        rom[151][19] = 16'hFFFE;
        rom[151][20] = 16'hFFE9;
        rom[151][21] = 16'hFFFA;
        rom[151][22] = 16'h000B;
        rom[151][23] = 16'hFFE0;
        rom[151][24] = 16'h0014;
        rom[151][25] = 16'hFFF4;
        rom[151][26] = 16'hFFFC;
        rom[151][27] = 16'hFFFA;
        rom[151][28] = 16'hFFF4;
        rom[151][29] = 16'hFFFE;
        rom[151][30] = 16'h0015;
        rom[151][31] = 16'h0002;
        rom[151][32] = 16'hFF9E;
        rom[151][33] = 16'h0001;
        rom[151][34] = 16'h001C;
        rom[151][35] = 16'h0015;
        rom[151][36] = 16'h0000;
        rom[151][37] = 16'h0012;
        rom[151][38] = 16'hFFE2;
        rom[151][39] = 16'h001A;
        rom[151][40] = 16'h000F;
        rom[151][41] = 16'hFFE6;
        rom[151][42] = 16'hFFF3;
        rom[151][43] = 16'hFFFA;
        rom[151][44] = 16'h0023;
        rom[151][45] = 16'hFFFA;
        rom[151][46] = 16'hFFE3;
        rom[151][47] = 16'h000D;
        rom[151][48] = 16'hFFF9;
        rom[151][49] = 16'h002D;
        rom[151][50] = 16'hFFDD;
        rom[151][51] = 16'h001D;
        rom[151][52] = 16'hFFB4;
        rom[151][53] = 16'hFFCE;
        rom[151][54] = 16'hFFDF;
        rom[151][55] = 16'h0002;
        rom[151][56] = 16'hFFE5;
        rom[151][57] = 16'hFFF1;
        rom[151][58] = 16'hFFF9;
        rom[151][59] = 16'hFFD5;
        rom[151][60] = 16'h0015;
        rom[151][61] = 16'hFFF7;
        rom[151][62] = 16'h000A;
        rom[151][63] = 16'hFFFE;
        rom[151][64] = 16'h000F;
        rom[151][65] = 16'hFFF9;
        rom[151][66] = 16'hFFE8;
        rom[151][67] = 16'h0012;
        rom[151][68] = 16'h002A;
        rom[151][69] = 16'h0015;
        rom[151][70] = 16'hFFF0;
        rom[151][71] = 16'hFFDA;
        rom[151][72] = 16'h0006;
        rom[151][73] = 16'h000B;
        rom[151][74] = 16'h0002;
        rom[151][75] = 16'h000C;
        rom[151][76] = 16'hFFCA;
        rom[151][77] = 16'hFFF3;
        rom[151][78] = 16'hFFFD;
        rom[151][79] = 16'h0003;
        rom[151][80] = 16'h0012;
        rom[151][81] = 16'hFFDC;
        rom[151][82] = 16'hFFB9;
        rom[151][83] = 16'h0002;
        rom[151][84] = 16'hFFDA;
        rom[151][85] = 16'hFFBF;
        rom[151][86] = 16'h0012;
        rom[151][87] = 16'h0005;
        rom[151][88] = 16'h000C;
        rom[151][89] = 16'hFFFD;
        rom[151][90] = 16'hFFF9;
        rom[151][91] = 16'hFFF3;
        rom[151][92] = 16'hFFF3;
        rom[151][93] = 16'h001B;
        rom[151][94] = 16'hFFBB;
        rom[151][95] = 16'h000D;
        rom[151][96] = 16'h000F;
        rom[151][97] = 16'hFFF1;
        rom[151][98] = 16'h0017;
        rom[151][99] = 16'h0002;
        rom[151][100] = 16'h001B;
        rom[151][101] = 16'hFFC9;
        rom[151][102] = 16'hFFEE;
        rom[151][103] = 16'h0027;
        rom[151][104] = 16'h0002;
        rom[151][105] = 16'hFFF3;
        rom[151][106] = 16'hFFC3;
        rom[151][107] = 16'h001A;
        rom[151][108] = 16'hFFEA;
        rom[151][109] = 16'h002B;
        rom[151][110] = 16'hFFDC;
        rom[151][111] = 16'h0002;
        rom[151][112] = 16'hFFC3;
        rom[151][113] = 16'hFFDE;
        rom[151][114] = 16'hFFFE;
        rom[151][115] = 16'h0004;
        rom[151][116] = 16'hFFEA;
        rom[151][117] = 16'hFFF9;
        rom[151][118] = 16'hFFC8;
        rom[151][119] = 16'hFFFC;
        rom[151][120] = 16'h000A;
        rom[151][121] = 16'h0032;
        rom[151][122] = 16'hFFD2;
        rom[151][123] = 16'hFFF0;
        rom[151][124] = 16'hFF98;
        rom[151][125] = 16'h0016;
        rom[151][126] = 16'h0011;
        rom[151][127] = 16'h0011;
        rom[152][0] = 16'h0016;
        rom[152][1] = 16'hFFF2;
        rom[152][2] = 16'h0008;
        rom[152][3] = 16'h000D;
        rom[152][4] = 16'hFFE5;
        rom[152][5] = 16'hFFE5;
        rom[152][6] = 16'h0014;
        rom[152][7] = 16'hFFF2;
        rom[152][8] = 16'h0011;
        rom[152][9] = 16'hFFDC;
        rom[152][10] = 16'h0025;
        rom[152][11] = 16'hFFEC;
        rom[152][12] = 16'hFFF6;
        rom[152][13] = 16'hFFF3;
        rom[152][14] = 16'hFFDB;
        rom[152][15] = 16'hFFED;
        rom[152][16] = 16'h0039;
        rom[152][17] = 16'h0019;
        rom[152][18] = 16'hFFE0;
        rom[152][19] = 16'h0019;
        rom[152][20] = 16'hFFBD;
        rom[152][21] = 16'h0000;
        rom[152][22] = 16'h0004;
        rom[152][23] = 16'hFFD5;
        rom[152][24] = 16'hFFFE;
        rom[152][25] = 16'hFFD3;
        rom[152][26] = 16'hFFF9;
        rom[152][27] = 16'hFFC9;
        rom[152][28] = 16'hFFFE;
        rom[152][29] = 16'h000F;
        rom[152][30] = 16'h0002;
        rom[152][31] = 16'h0019;
        rom[152][32] = 16'hFFD1;
        rom[152][33] = 16'hFFDE;
        rom[152][34] = 16'hFFF3;
        rom[152][35] = 16'h000D;
        rom[152][36] = 16'hFFE7;
        rom[152][37] = 16'h0013;
        rom[152][38] = 16'hFFF2;
        rom[152][39] = 16'h0015;
        rom[152][40] = 16'hFFFC;
        rom[152][41] = 16'hFFD9;
        rom[152][42] = 16'h0016;
        rom[152][43] = 16'hFFC1;
        rom[152][44] = 16'h002B;
        rom[152][45] = 16'h0009;
        rom[152][46] = 16'hFFC7;
        rom[152][47] = 16'hFFF7;
        rom[152][48] = 16'h0003;
        rom[152][49] = 16'h0005;
        rom[152][50] = 16'h000E;
        rom[152][51] = 16'h0004;
        rom[152][52] = 16'hFFF3;
        rom[152][53] = 16'hFFD8;
        rom[152][54] = 16'hFFD0;
        rom[152][55] = 16'h0002;
        rom[152][56] = 16'hFFFB;
        rom[152][57] = 16'hFFEA;
        rom[152][58] = 16'hFFE9;
        rom[152][59] = 16'hFFED;
        rom[152][60] = 16'h0001;
        rom[152][61] = 16'hFFE7;
        rom[152][62] = 16'h0000;
        rom[152][63] = 16'hFFED;
        rom[152][64] = 16'h000F;
        rom[152][65] = 16'hFFEA;
        rom[152][66] = 16'hFFFD;
        rom[152][67] = 16'hFFDB;
        rom[152][68] = 16'h000E;
        rom[152][69] = 16'h0024;
        rom[152][70] = 16'h000C;
        rom[152][71] = 16'h0009;
        rom[152][72] = 16'hFFE0;
        rom[152][73] = 16'hFFFD;
        rom[152][74] = 16'hFFED;
        rom[152][75] = 16'hFFAB;
        rom[152][76] = 16'hFFE9;
        rom[152][77] = 16'h0002;
        rom[152][78] = 16'h0017;
        rom[152][79] = 16'h001B;
        rom[152][80] = 16'hFFF1;
        rom[152][81] = 16'hFF98;
        rom[152][82] = 16'h0002;
        rom[152][83] = 16'hFFF2;
        rom[152][84] = 16'hFFD3;
        rom[152][85] = 16'hFFE1;
        rom[152][86] = 16'h001D;
        rom[152][87] = 16'hFFF8;
        rom[152][88] = 16'h0006;
        rom[152][89] = 16'hFFEF;
        rom[152][90] = 16'hFFC5;
        rom[152][91] = 16'h0021;
        rom[152][92] = 16'hFFF0;
        rom[152][93] = 16'h002A;
        rom[152][94] = 16'h0001;
        rom[152][95] = 16'hFFFF;
        rom[152][96] = 16'h002E;
        rom[152][97] = 16'h000C;
        rom[152][98] = 16'h001F;
        rom[152][99] = 16'hFFBA;
        rom[152][100] = 16'h003A;
        rom[152][101] = 16'hFFF3;
        rom[152][102] = 16'h000A;
        rom[152][103] = 16'h001A;
        rom[152][104] = 16'hFFEC;
        rom[152][105] = 16'h0007;
        rom[152][106] = 16'h001E;
        rom[152][107] = 16'hFFEF;
        rom[152][108] = 16'hFFE6;
        rom[152][109] = 16'h000C;
        rom[152][110] = 16'hFFE6;
        rom[152][111] = 16'h0012;
        rom[152][112] = 16'hFFEF;
        rom[152][113] = 16'hFFF9;
        rom[152][114] = 16'hFFDF;
        rom[152][115] = 16'h0001;
        rom[152][116] = 16'hFFE5;
        rom[152][117] = 16'h0008;
        rom[152][118] = 16'hFFEF;
        rom[152][119] = 16'hFFD2;
        rom[152][120] = 16'hFFC6;
        rom[152][121] = 16'h001F;
        rom[152][122] = 16'hFFE5;
        rom[152][123] = 16'hFFEB;
        rom[152][124] = 16'hFFEE;
        rom[152][125] = 16'hFFF6;
        rom[152][126] = 16'h0034;
        rom[152][127] = 16'h0003;
        rom[153][0] = 16'h0003;
        rom[153][1] = 16'hFFF6;
        rom[153][2] = 16'hFFD0;
        rom[153][3] = 16'h000A;
        rom[153][4] = 16'hFFF0;
        rom[153][5] = 16'h0014;
        rom[153][6] = 16'h0004;
        rom[153][7] = 16'h0009;
        rom[153][8] = 16'hFFE1;
        rom[153][9] = 16'h0017;
        rom[153][10] = 16'h0018;
        rom[153][11] = 16'h004B;
        rom[153][12] = 16'h0008;
        rom[153][13] = 16'h001F;
        rom[153][14] = 16'h0001;
        rom[153][15] = 16'hFFE9;
        rom[153][16] = 16'h0028;
        rom[153][17] = 16'hFFF9;
        rom[153][18] = 16'h0011;
        rom[153][19] = 16'h000A;
        rom[153][20] = 16'hFFEE;
        rom[153][21] = 16'hFFC8;
        rom[153][22] = 16'h0007;
        rom[153][23] = 16'h000D;
        rom[153][24] = 16'hFFE9;
        rom[153][25] = 16'hFFEA;
        rom[153][26] = 16'hFFDE;
        rom[153][27] = 16'hFFC9;
        rom[153][28] = 16'hFFEC;
        rom[153][29] = 16'hFFEF;
        rom[153][30] = 16'hFFFC;
        rom[153][31] = 16'hFFF6;
        rom[153][32] = 16'h0017;
        rom[153][33] = 16'h0009;
        rom[153][34] = 16'hFFF4;
        rom[153][35] = 16'hFFFB;
        rom[153][36] = 16'h001F;
        rom[153][37] = 16'hFFF4;
        rom[153][38] = 16'h002E;
        rom[153][39] = 16'hFFCF;
        rom[153][40] = 16'h0007;
        rom[153][41] = 16'hFFDD;
        rom[153][42] = 16'h000B;
        rom[153][43] = 16'h0022;
        rom[153][44] = 16'hFFFC;
        rom[153][45] = 16'h0004;
        rom[153][46] = 16'h0028;
        rom[153][47] = 16'hFFF8;
        rom[153][48] = 16'h003D;
        rom[153][49] = 16'hFFE7;
        rom[153][50] = 16'h002A;
        rom[153][51] = 16'h0011;
        rom[153][52] = 16'hFFEF;
        rom[153][53] = 16'h0009;
        rom[153][54] = 16'hFFEB;
        rom[153][55] = 16'hFFFE;
        rom[153][56] = 16'hFFE2;
        rom[153][57] = 16'h0011;
        rom[153][58] = 16'hFFF4;
        rom[153][59] = 16'h0013;
        rom[153][60] = 16'hFFF5;
        rom[153][61] = 16'h0001;
        rom[153][62] = 16'hFFD3;
        rom[153][63] = 16'h0003;
        rom[153][64] = 16'hFFD2;
        rom[153][65] = 16'h0024;
        rom[153][66] = 16'hFFBA;
        rom[153][67] = 16'hFFCE;
        rom[153][68] = 16'hFFFD;
        rom[153][69] = 16'hFFE6;
        rom[153][70] = 16'hFFCE;
        rom[153][71] = 16'hFFD9;
        rom[153][72] = 16'hFFD5;
        rom[153][73] = 16'hFFC5;
        rom[153][74] = 16'h0007;
        rom[153][75] = 16'hFFEA;
        rom[153][76] = 16'hFFDC;
        rom[153][77] = 16'hFFFB;
        rom[153][78] = 16'hFFEE;
        rom[153][79] = 16'hFFD4;
        rom[153][80] = 16'hFFF5;
        rom[153][81] = 16'hFFFE;
        rom[153][82] = 16'hFFF9;
        rom[153][83] = 16'hFFEC;
        rom[153][84] = 16'h0030;
        rom[153][85] = 16'h002E;
        rom[153][86] = 16'hFFEF;
        rom[153][87] = 16'h000B;
        rom[153][88] = 16'hFFF8;
        rom[153][89] = 16'hFFEF;
        rom[153][90] = 16'h0016;
        rom[153][91] = 16'h0009;
        rom[153][92] = 16'hFFFE;
        rom[153][93] = 16'hFFCB;
        rom[153][94] = 16'hFFEA;
        rom[153][95] = 16'h0027;
        rom[153][96] = 16'h0005;
        rom[153][97] = 16'hFFAF;
        rom[153][98] = 16'hFFE3;
        rom[153][99] = 16'h002B;
        rom[153][100] = 16'hFFEC;
        rom[153][101] = 16'hFFF9;
        rom[153][102] = 16'h000C;
        rom[153][103] = 16'h000B;
        rom[153][104] = 16'hFFEF;
        rom[153][105] = 16'h001C;
        rom[153][106] = 16'hFFF8;
        rom[153][107] = 16'hFFE5;
        rom[153][108] = 16'hFFE6;
        rom[153][109] = 16'hFFED;
        rom[153][110] = 16'h001C;
        rom[153][111] = 16'hFFDE;
        rom[153][112] = 16'hFFCF;
        rom[153][113] = 16'hFFFB;
        rom[153][114] = 16'hFFCD;
        rom[153][115] = 16'hFFFB;
        rom[153][116] = 16'h001F;
        rom[153][117] = 16'hFFFF;
        rom[153][118] = 16'hFFF5;
        rom[153][119] = 16'hFFF8;
        rom[153][120] = 16'h0029;
        rom[153][121] = 16'h0031;
        rom[153][122] = 16'hFFF4;
        rom[153][123] = 16'h002A;
        rom[153][124] = 16'hFFF1;
        rom[153][125] = 16'hFFF1;
        rom[153][126] = 16'hFFF4;
        rom[153][127] = 16'h0004;
        rom[154][0] = 16'hFFDE;
        rom[154][1] = 16'h0031;
        rom[154][2] = 16'h0015;
        rom[154][3] = 16'h002D;
        rom[154][4] = 16'hFFC1;
        rom[154][5] = 16'h001F;
        rom[154][6] = 16'h0007;
        rom[154][7] = 16'h0006;
        rom[154][8] = 16'h000E;
        rom[154][9] = 16'hFFE1;
        rom[154][10] = 16'hFFD5;
        rom[154][11] = 16'h001F;
        rom[154][12] = 16'hFFCA;
        rom[154][13] = 16'hFFF9;
        rom[154][14] = 16'hFFC3;
        rom[154][15] = 16'hFFE1;
        rom[154][16] = 16'h0007;
        rom[154][17] = 16'hFFDE;
        rom[154][18] = 16'hFFE2;
        rom[154][19] = 16'h000C;
        rom[154][20] = 16'h0024;
        rom[154][21] = 16'h0002;
        rom[154][22] = 16'hFFDC;
        rom[154][23] = 16'hFFE4;
        rom[154][24] = 16'h0002;
        rom[154][25] = 16'h0010;
        rom[154][26] = 16'h0009;
        rom[154][27] = 16'hFFF4;
        rom[154][28] = 16'hFFC2;
        rom[154][29] = 16'hFFF4;
        rom[154][30] = 16'hFFFA;
        rom[154][31] = 16'hFFEC;
        rom[154][32] = 16'hFFFD;
        rom[154][33] = 16'hFFB8;
        rom[154][34] = 16'h001F;
        rom[154][35] = 16'hFFC2;
        rom[154][36] = 16'h001C;
        rom[154][37] = 16'hFFD1;
        rom[154][38] = 16'hFFEB;
        rom[154][39] = 16'h000D;
        rom[154][40] = 16'h001E;
        rom[154][41] = 16'hFFE8;
        rom[154][42] = 16'hFFC6;
        rom[154][43] = 16'h0028;
        rom[154][44] = 16'hFFF9;
        rom[154][45] = 16'hFFBF;
        rom[154][46] = 16'h0018;
        rom[154][47] = 16'h0034;
        rom[154][48] = 16'h001B;
        rom[154][49] = 16'hFFE9;
        rom[154][50] = 16'h001E;
        rom[154][51] = 16'h0004;
        rom[154][52] = 16'hFFEF;
        rom[154][53] = 16'h0019;
        rom[154][54] = 16'h000F;
        rom[154][55] = 16'h002B;
        rom[154][56] = 16'hFFE5;
        rom[154][57] = 16'hFFBE;
        rom[154][58] = 16'hFFF7;
        rom[154][59] = 16'hFFF9;
        rom[154][60] = 16'h0008;
        rom[154][61] = 16'hFFFE;
        rom[154][62] = 16'h002B;
        rom[154][63] = 16'h0025;
        rom[154][64] = 16'hFFF9;
        rom[154][65] = 16'hFFF5;
        rom[154][66] = 16'hFFF4;
        rom[154][67] = 16'h001B;
        rom[154][68] = 16'h000A;
        rom[154][69] = 16'h0012;
        rom[154][70] = 16'h000A;
        rom[154][71] = 16'hFFD9;
        rom[154][72] = 16'hFFE0;
        rom[154][73] = 16'hFFDB;
        rom[154][74] = 16'h000E;
        rom[154][75] = 16'hFFA7;
        rom[154][76] = 16'h0007;
        rom[154][77] = 16'hFFD8;
        rom[154][78] = 16'h0011;
        rom[154][79] = 16'hFFFE;
        rom[154][80] = 16'h0023;
        rom[154][81] = 16'hFFE0;
        rom[154][82] = 16'h002E;
        rom[154][83] = 16'h0017;
        rom[154][84] = 16'hFFCC;
        rom[154][85] = 16'h0000;
        rom[154][86] = 16'h000D;
        rom[154][87] = 16'h0009;
        rom[154][88] = 16'h0037;
        rom[154][89] = 16'hFFC4;
        rom[154][90] = 16'h000F;
        rom[154][91] = 16'h0017;
        rom[154][92] = 16'hFFF3;
        rom[154][93] = 16'h0006;
        rom[154][94] = 16'hFFE8;
        rom[154][95] = 16'hFFBA;
        rom[154][96] = 16'h000F;
        rom[154][97] = 16'h0022;
        rom[154][98] = 16'h000F;
        rom[154][99] = 16'hFFFB;
        rom[154][100] = 16'hFFED;
        rom[154][101] = 16'h0018;
        rom[154][102] = 16'h0012;
        rom[154][103] = 16'hFFFE;
        rom[154][104] = 16'hFFE5;
        rom[154][105] = 16'hFFE7;
        rom[154][106] = 16'h0026;
        rom[154][107] = 16'hFFD2;
        rom[154][108] = 16'hFFEA;
        rom[154][109] = 16'hFFE2;
        rom[154][110] = 16'hFFF9;
        rom[154][111] = 16'h0008;
        rom[154][112] = 16'h0026;
        rom[154][113] = 16'hFFFE;
        rom[154][114] = 16'hFFDD;
        rom[154][115] = 16'h001B;
        rom[154][116] = 16'hFFE7;
        rom[154][117] = 16'hFFF4;
        rom[154][118] = 16'h0007;
        rom[154][119] = 16'hFFD6;
        rom[154][120] = 16'h0023;
        rom[154][121] = 16'h001D;
        rom[154][122] = 16'h0012;
        rom[154][123] = 16'hFFDC;
        rom[154][124] = 16'hFFF0;
        rom[154][125] = 16'hFFF4;
        rom[154][126] = 16'hFFFC;
        rom[154][127] = 16'h0009;
        rom[155][0] = 16'h0011;
        rom[155][1] = 16'h0023;
        rom[155][2] = 16'hFFD8;
        rom[155][3] = 16'h0028;
        rom[155][4] = 16'h000B;
        rom[155][5] = 16'h000C;
        rom[155][6] = 16'h0010;
        rom[155][7] = 16'hFFFA;
        rom[155][8] = 16'hFFD2;
        rom[155][9] = 16'hFFDC;
        rom[155][10] = 16'h000A;
        rom[155][11] = 16'hFFD1;
        rom[155][12] = 16'h0014;
        rom[155][13] = 16'h0009;
        rom[155][14] = 16'hFFEF;
        rom[155][15] = 16'hFFCD;
        rom[155][16] = 16'h0032;
        rom[155][17] = 16'hFFDF;
        rom[155][18] = 16'hFFF2;
        rom[155][19] = 16'hFFFE;
        rom[155][20] = 16'hFFE0;
        rom[155][21] = 16'hFFB9;
        rom[155][22] = 16'hFFFE;
        rom[155][23] = 16'h0027;
        rom[155][24] = 16'hFFDE;
        rom[155][25] = 16'h0016;
        rom[155][26] = 16'h0023;
        rom[155][27] = 16'hFFE9;
        rom[155][28] = 16'hFFDD;
        rom[155][29] = 16'hFFF4;
        rom[155][30] = 16'hFFEA;
        rom[155][31] = 16'hFFF9;
        rom[155][32] = 16'hFFE1;
        rom[155][33] = 16'hFFDB;
        rom[155][34] = 16'hFFF7;
        rom[155][35] = 16'hFFBD;
        rom[155][36] = 16'h0016;
        rom[155][37] = 16'hFFEC;
        rom[155][38] = 16'hFFE0;
        rom[155][39] = 16'hFFE6;
        rom[155][40] = 16'h003E;
        rom[155][41] = 16'h0001;
        rom[155][42] = 16'h0016;
        rom[155][43] = 16'hFFD9;
        rom[155][44] = 16'hFFF8;
        rom[155][45] = 16'hFFBA;
        rom[155][46] = 16'h003A;
        rom[155][47] = 16'h0008;
        rom[155][48] = 16'h0010;
        rom[155][49] = 16'h0036;
        rom[155][50] = 16'hFFE7;
        rom[155][51] = 16'hFFF3;
        rom[155][52] = 16'hFFD5;
        rom[155][53] = 16'hFFF1;
        rom[155][54] = 16'hFFF0;
        rom[155][55] = 16'hFFE9;
        rom[155][56] = 16'hFFE2;
        rom[155][57] = 16'h000A;
        rom[155][58] = 16'h0016;
        rom[155][59] = 16'hFFCE;
        rom[155][60] = 16'hFFE5;
        rom[155][61] = 16'hFFE3;
        rom[155][62] = 16'h0002;
        rom[155][63] = 16'hFFF3;
        rom[155][64] = 16'hFFFA;
        rom[155][65] = 16'hFFE2;
        rom[155][66] = 16'h0006;
        rom[155][67] = 16'h001B;
        rom[155][68] = 16'h0008;
        rom[155][69] = 16'h0007;
        rom[155][70] = 16'hFFE4;
        rom[155][71] = 16'hFFEF;
        rom[155][72] = 16'h0009;
        rom[155][73] = 16'h0013;
        rom[155][74] = 16'h0005;
        rom[155][75] = 16'hFFC5;
        rom[155][76] = 16'hFFD8;
        rom[155][77] = 16'h0002;
        rom[155][78] = 16'h0007;
        rom[155][79] = 16'h0001;
        rom[155][80] = 16'hFFF6;
        rom[155][81] = 16'h000B;
        rom[155][82] = 16'h0024;
        rom[155][83] = 16'h0005;
        rom[155][84] = 16'hFFE9;
        rom[155][85] = 16'hFFFE;
        rom[155][86] = 16'h001C;
        rom[155][87] = 16'hFFEB;
        rom[155][88] = 16'hFFEB;
        rom[155][89] = 16'hFFDF;
        rom[155][90] = 16'h0000;
        rom[155][91] = 16'h002F;
        rom[155][92] = 16'h0008;
        rom[155][93] = 16'hFFE4;
        rom[155][94] = 16'hFFF4;
        rom[155][95] = 16'h001C;
        rom[155][96] = 16'hFFF7;
        rom[155][97] = 16'hFFEB;
        rom[155][98] = 16'h0022;
        rom[155][99] = 16'h0015;
        rom[155][100] = 16'h0007;
        rom[155][101] = 16'h001B;
        rom[155][102] = 16'h002A;
        rom[155][103] = 16'hFFFD;
        rom[155][104] = 16'h0026;
        rom[155][105] = 16'hFFE4;
        rom[155][106] = 16'h0004;
        rom[155][107] = 16'hFFBF;
        rom[155][108] = 16'h0002;
        rom[155][109] = 16'hFFE5;
        rom[155][110] = 16'hFFE2;
        rom[155][111] = 16'hFFFE;
        rom[155][112] = 16'h001B;
        rom[155][113] = 16'h002C;
        rom[155][114] = 16'h0005;
        rom[155][115] = 16'hFFEF;
        rom[155][116] = 16'hFFC4;
        rom[155][117] = 16'h000E;
        rom[155][118] = 16'hFFE3;
        rom[155][119] = 16'hFFC3;
        rom[155][120] = 16'h0002;
        rom[155][121] = 16'h0015;
        rom[155][122] = 16'hFFD2;
        rom[155][123] = 16'h0018;
        rom[155][124] = 16'h0007;
        rom[155][125] = 16'h0024;
        rom[155][126] = 16'hFFE6;
        rom[155][127] = 16'hFFEA;
        rom[156][0] = 16'h0011;
        rom[156][1] = 16'hFFF7;
        rom[156][2] = 16'hFFC3;
        rom[156][3] = 16'hFFE7;
        rom[156][4] = 16'hFFE9;
        rom[156][5] = 16'hFFC1;
        rom[156][6] = 16'h000F;
        rom[156][7] = 16'h001B;
        rom[156][8] = 16'h0033;
        rom[156][9] = 16'hFFF2;
        rom[156][10] = 16'h001A;
        rom[156][11] = 16'h0011;
        rom[156][12] = 16'hFFF1;
        rom[156][13] = 16'h000D;
        rom[156][14] = 16'hFFDD;
        rom[156][15] = 16'hFFE7;
        rom[156][16] = 16'h0024;
        rom[156][17] = 16'h0014;
        rom[156][18] = 16'h001E;
        rom[156][19] = 16'hFFE7;
        rom[156][20] = 16'hFFCE;
        rom[156][21] = 16'h0018;
        rom[156][22] = 16'h0014;
        rom[156][23] = 16'h0015;
        rom[156][24] = 16'h001B;
        rom[156][25] = 16'hFFB5;
        rom[156][26] = 16'hFFFB;
        rom[156][27] = 16'hFFCA;
        rom[156][28] = 16'h0023;
        rom[156][29] = 16'h0019;
        rom[156][30] = 16'hFFF3;
        rom[156][31] = 16'h0006;
        rom[156][32] = 16'hFFEA;
        rom[156][33] = 16'h0044;
        rom[156][34] = 16'hFFF5;
        rom[156][35] = 16'h0013;
        rom[156][36] = 16'h0001;
        rom[156][37] = 16'hFFFE;
        rom[156][38] = 16'h0006;
        rom[156][39] = 16'h0022;
        rom[156][40] = 16'h000E;
        rom[156][41] = 16'h0021;
        rom[156][42] = 16'hFFDF;
        rom[156][43] = 16'hFFD9;
        rom[156][44] = 16'h001F;
        rom[156][45] = 16'hFFEE;
        rom[156][46] = 16'hFFFF;
        rom[156][47] = 16'hFFEF;
        rom[156][48] = 16'hFFE5;
        rom[156][49] = 16'hFFFB;
        rom[156][50] = 16'hFFD2;
        rom[156][51] = 16'hFFE1;
        rom[156][52] = 16'hFFE5;
        rom[156][53] = 16'hFFF2;
        rom[156][54] = 16'hFFCE;
        rom[156][55] = 16'hFFD2;
        rom[156][56] = 16'hFFF8;
        rom[156][57] = 16'h000C;
        rom[156][58] = 16'h0000;
        rom[156][59] = 16'hFFC9;
        rom[156][60] = 16'h0009;
        rom[156][61] = 16'hFFFF;
        rom[156][62] = 16'hFFF9;
        rom[156][63] = 16'hFFE4;
        rom[156][64] = 16'hFFFA;
        rom[156][65] = 16'h000E;
        rom[156][66] = 16'hFFB6;
        rom[156][67] = 16'hFFD7;
        rom[156][68] = 16'h0041;
        rom[156][69] = 16'hFFE7;
        rom[156][70] = 16'h000D;
        rom[156][71] = 16'hFFD3;
        rom[156][72] = 16'h000B;
        rom[156][73] = 16'hFFE0;
        rom[156][74] = 16'h000D;
        rom[156][75] = 16'h0007;
        rom[156][76] = 16'hFFDE;
        rom[156][77] = 16'hFFED;
        rom[156][78] = 16'h000C;
        rom[156][79] = 16'hFFC0;
        rom[156][80] = 16'hFFFE;
        rom[156][81] = 16'hFFDA;
        rom[156][82] = 16'hFFDC;
        rom[156][83] = 16'h0004;
        rom[156][84] = 16'h0013;
        rom[156][85] = 16'hFFEB;
        rom[156][86] = 16'h0023;
        rom[156][87] = 16'hFFF4;
        rom[156][88] = 16'hFFF4;
        rom[156][89] = 16'h0011;
        rom[156][90] = 16'hFFD4;
        rom[156][91] = 16'h0011;
        rom[156][92] = 16'h002C;
        rom[156][93] = 16'h001A;
        rom[156][94] = 16'h0033;
        rom[156][95] = 16'h001A;
        rom[156][96] = 16'h0012;
        rom[156][97] = 16'h0029;
        rom[156][98] = 16'h001B;
        rom[156][99] = 16'h002A;
        rom[156][100] = 16'hFFFD;
        rom[156][101] = 16'hFFDC;
        rom[156][102] = 16'hFFEA;
        rom[156][103] = 16'hFFE5;
        rom[156][104] = 16'hFFE6;
        rom[156][105] = 16'h000B;
        rom[156][106] = 16'hFFBB;
        rom[156][107] = 16'hFFE2;
        rom[156][108] = 16'h0016;
        rom[156][109] = 16'h0018;
        rom[156][110] = 16'h000C;
        rom[156][111] = 16'hFFF1;
        rom[156][112] = 16'hFFF9;
        rom[156][113] = 16'hFFF7;
        rom[156][114] = 16'hFFFF;
        rom[156][115] = 16'hFFF0;
        rom[156][116] = 16'h002E;
        rom[156][117] = 16'h0017;
        rom[156][118] = 16'hFFC8;
        rom[156][119] = 16'hFFD5;
        rom[156][120] = 16'h0007;
        rom[156][121] = 16'h0015;
        rom[156][122] = 16'h000B;
        rom[156][123] = 16'h0016;
        rom[156][124] = 16'hFFF4;
        rom[156][125] = 16'hFFD0;
        rom[156][126] = 16'hFFE6;
        rom[156][127] = 16'h000F;
        rom[157][0] = 16'h0007;
        rom[157][1] = 16'h001A;
        rom[157][2] = 16'h0002;
        rom[157][3] = 16'hFFDA;
        rom[157][4] = 16'hFFEA;
        rom[157][5] = 16'hFFC8;
        rom[157][6] = 16'hFFE7;
        rom[157][7] = 16'h0013;
        rom[157][8] = 16'hFFF6;
        rom[157][9] = 16'h000B;
        rom[157][10] = 16'h0002;
        rom[157][11] = 16'hFFF1;
        rom[157][12] = 16'hFFE5;
        rom[157][13] = 16'h0008;
        rom[157][14] = 16'h0006;
        rom[157][15] = 16'h002E;
        rom[157][16] = 16'hFFEF;
        rom[157][17] = 16'hFFFF;
        rom[157][18] = 16'hFFFE;
        rom[157][19] = 16'h000E;
        rom[157][20] = 16'h0002;
        rom[157][21] = 16'h0016;
        rom[157][22] = 16'h0012;
        rom[157][23] = 16'h001A;
        rom[157][24] = 16'h0002;
        rom[157][25] = 16'hFFB2;
        rom[157][26] = 16'hFFE5;
        rom[157][27] = 16'hFFDC;
        rom[157][28] = 16'hFFEE;
        rom[157][29] = 16'h000C;
        rom[157][30] = 16'hFFD8;
        rom[157][31] = 16'h003B;
        rom[157][32] = 16'hFFF3;
        rom[157][33] = 16'hFFFF;
        rom[157][34] = 16'h000C;
        rom[157][35] = 16'hFFF8;
        rom[157][36] = 16'hFFF0;
        rom[157][37] = 16'hFFF9;
        rom[157][38] = 16'h000C;
        rom[157][39] = 16'h003D;
        rom[157][40] = 16'hFFD7;
        rom[157][41] = 16'h0028;
        rom[157][42] = 16'h0021;
        rom[157][43] = 16'hFFFB;
        rom[157][44] = 16'h0030;
        rom[157][45] = 16'hFFB1;
        rom[157][46] = 16'hFFF9;
        rom[157][47] = 16'hFFE4;
        rom[157][48] = 16'hFFDE;
        rom[157][49] = 16'hFFE2;
        rom[157][50] = 16'hFFEC;
        rom[157][51] = 16'hFFEA;
        rom[157][52] = 16'h001E;
        rom[157][53] = 16'hFFE5;
        rom[157][54] = 16'hFFC6;
        rom[157][55] = 16'h001F;
        rom[157][56] = 16'h0009;
        rom[157][57] = 16'h0025;
        rom[157][58] = 16'h0002;
        rom[157][59] = 16'hFFF8;
        rom[157][60] = 16'h0002;
        rom[157][61] = 16'hFFE1;
        rom[157][62] = 16'hFFC8;
        rom[157][63] = 16'hFFB8;
        rom[157][64] = 16'h001A;
        rom[157][65] = 16'h001A;
        rom[157][66] = 16'hFFDE;
        rom[157][67] = 16'hFFE1;
        rom[157][68] = 16'hFFED;
        rom[157][69] = 16'h001F;
        rom[157][70] = 16'h0016;
        rom[157][71] = 16'h001D;
        rom[157][72] = 16'hFFEB;
        rom[157][73] = 16'hFFE5;
        rom[157][74] = 16'h0026;
        rom[157][75] = 16'hFFEF;
        rom[157][76] = 16'h001F;
        rom[157][77] = 16'hFFFA;
        rom[157][78] = 16'h0029;
        rom[157][79] = 16'hFFE1;
        rom[157][80] = 16'h0018;
        rom[157][81] = 16'hFFBF;
        rom[157][82] = 16'hFFDC;
        rom[157][83] = 16'hFFF1;
        rom[157][84] = 16'h000E;
        rom[157][85] = 16'hFFEC;
        rom[157][86] = 16'hFFF2;
        rom[157][87] = 16'hFFF2;
        rom[157][88] = 16'hFFFA;
        rom[157][89] = 16'hFFAD;
        rom[157][90] = 16'hFFD0;
        rom[157][91] = 16'h0001;
        rom[157][92] = 16'hFFDC;
        rom[157][93] = 16'hFFE5;
        rom[157][94] = 16'h0011;
        rom[157][95] = 16'h0015;
        rom[157][96] = 16'hFFE7;
        rom[157][97] = 16'hFFCD;
        rom[157][98] = 16'hFFCE;
        rom[157][99] = 16'hFFE6;
        rom[157][100] = 16'h002C;
        rom[157][101] = 16'h0012;
        rom[157][102] = 16'hFFF4;
        rom[157][103] = 16'h001F;
        rom[157][104] = 16'hFFEA;
        rom[157][105] = 16'h000C;
        rom[157][106] = 16'hFFEE;
        rom[157][107] = 16'hFFF4;
        rom[157][108] = 16'hFFF2;
        rom[157][109] = 16'h0006;
        rom[157][110] = 16'hFFE9;
        rom[157][111] = 16'hFFCE;
        rom[157][112] = 16'h0014;
        rom[157][113] = 16'hFFF4;
        rom[157][114] = 16'h0007;
        rom[157][115] = 16'hFFF8;
        rom[157][116] = 16'hFFFA;
        rom[157][117] = 16'h001E;
        rom[157][118] = 16'hFFB4;
        rom[157][119] = 16'h0004;
        rom[157][120] = 16'hFFE7;
        rom[157][121] = 16'h0011;
        rom[157][122] = 16'h000C;
        rom[157][123] = 16'hFFF9;
        rom[157][124] = 16'hFFD2;
        rom[157][125] = 16'hFFDB;
        rom[157][126] = 16'h0003;
        rom[157][127] = 16'h001B;
        rom[158][0] = 16'h0001;
        rom[158][1] = 16'h001D;
        rom[158][2] = 16'hFFDC;
        rom[158][3] = 16'hFFD0;
        rom[158][4] = 16'hFFEC;
        rom[158][5] = 16'hFFE5;
        rom[158][6] = 16'hFFEA;
        rom[158][7] = 16'h000D;
        rom[158][8] = 16'h0011;
        rom[158][9] = 16'hFFF3;
        rom[158][10] = 16'h0026;
        rom[158][11] = 16'hFFF1;
        rom[158][12] = 16'h000D;
        rom[158][13] = 16'hFFDC;
        rom[158][14] = 16'h002A;
        rom[158][15] = 16'h000D;
        rom[158][16] = 16'hFFEF;
        rom[158][17] = 16'hFFE7;
        rom[158][18] = 16'h000D;
        rom[158][19] = 16'h0016;
        rom[158][20] = 16'h0006;
        rom[158][21] = 16'h0010;
        rom[158][22] = 16'hFFE2;
        rom[158][23] = 16'h0020;
        rom[158][24] = 16'h0011;
        rom[158][25] = 16'hFFE2;
        rom[158][26] = 16'h003F;
        rom[158][27] = 16'hFFAF;
        rom[158][28] = 16'hFFE7;
        rom[158][29] = 16'hFFFE;
        rom[158][30] = 16'h001B;
        rom[158][31] = 16'h0039;
        rom[158][32] = 16'h001F;
        rom[158][33] = 16'hFFFF;
        rom[158][34] = 16'hFFF7;
        rom[158][35] = 16'h0014;
        rom[158][36] = 16'h0012;
        rom[158][37] = 16'hFFE2;
        rom[158][38] = 16'hFFE5;
        rom[158][39] = 16'hFFEC;
        rom[158][40] = 16'hFFBF;
        rom[158][41] = 16'h001B;
        rom[158][42] = 16'hFFF4;
        rom[158][43] = 16'h000F;
        rom[158][44] = 16'hFFF8;
        rom[158][45] = 16'h002E;
        rom[158][46] = 16'h001B;
        rom[158][47] = 16'h0033;
        rom[158][48] = 16'hFFF9;
        rom[158][49] = 16'hFFEA;
        rom[158][50] = 16'hFFFE;
        rom[158][51] = 16'hFFDE;
        rom[158][52] = 16'hFFD1;
        rom[158][53] = 16'hFFCC;
        rom[158][54] = 16'hFFF9;
        rom[158][55] = 16'hFFC8;
        rom[158][56] = 16'hFFEF;
        rom[158][57] = 16'hFFD1;
        rom[158][58] = 16'h000B;
        rom[158][59] = 16'hFFF4;
        rom[158][60] = 16'h0013;
        rom[158][61] = 16'hFFFE;
        rom[158][62] = 16'h0003;
        rom[158][63] = 16'h0021;
        rom[158][64] = 16'hFFFE;
        rom[158][65] = 16'h0024;
        rom[158][66] = 16'hFFD4;
        rom[158][67] = 16'hFFEA;
        rom[158][68] = 16'hFFE2;
        rom[158][69] = 16'hFFF9;
        rom[158][70] = 16'h0030;
        rom[158][71] = 16'hFFCF;
        rom[158][72] = 16'h001E;
        rom[158][73] = 16'hFFF6;
        rom[158][74] = 16'h0026;
        rom[158][75] = 16'h0007;
        rom[158][76] = 16'hFFE1;
        rom[158][77] = 16'hFFDC;
        rom[158][78] = 16'h0040;
        rom[158][79] = 16'h002C;
        rom[158][80] = 16'hFFDE;
        rom[158][81] = 16'h002D;
        rom[158][82] = 16'h0012;
        rom[158][83] = 16'hFFFC;
        rom[158][84] = 16'h000C;
        rom[158][85] = 16'hFFD6;
        rom[158][86] = 16'hFFF2;
        rom[158][87] = 16'hFFCB;
        rom[158][88] = 16'hFFEC;
        rom[158][89] = 16'hFFFD;
        rom[158][90] = 16'h0014;
        rom[158][91] = 16'h0022;
        rom[158][92] = 16'h0019;
        rom[158][93] = 16'h0016;
        rom[158][94] = 16'hFFF6;
        rom[158][95] = 16'h0011;
        rom[158][96] = 16'h0005;
        rom[158][97] = 16'hFFEF;
        rom[158][98] = 16'h0009;
        rom[158][99] = 16'h0036;
        rom[158][100] = 16'hFFB5;
        rom[158][101] = 16'hFFF0;
        rom[158][102] = 16'hFFF0;
        rom[158][103] = 16'hFFD8;
        rom[158][104] = 16'hFFFF;
        rom[158][105] = 16'hFFE2;
        rom[158][106] = 16'hFFCB;
        rom[158][107] = 16'hFFF8;
        rom[158][108] = 16'hFFD1;
        rom[158][109] = 16'h0024;
        rom[158][110] = 16'hFFFE;
        rom[158][111] = 16'h002B;
        rom[158][112] = 16'hFFF9;
        rom[158][113] = 16'hFFFB;
        rom[158][114] = 16'hFFCF;
        rom[158][115] = 16'h0015;
        rom[158][116] = 16'h0007;
        rom[158][117] = 16'h0018;
        rom[158][118] = 16'h0024;
        rom[158][119] = 16'h0002;
        rom[158][120] = 16'hFFD6;
        rom[158][121] = 16'hFFFF;
        rom[158][122] = 16'hFFF7;
        rom[158][123] = 16'hFFF4;
        rom[158][124] = 16'hFFF5;
        rom[158][125] = 16'hFFFD;
        rom[158][126] = 16'hFFE8;
        rom[158][127] = 16'hFFFD;
        rom[159][0] = 16'hFFF8;
        rom[159][1] = 16'h0016;
        rom[159][2] = 16'hFFEC;
        rom[159][3] = 16'hFFFF;
        rom[159][4] = 16'hFFF3;
        rom[159][5] = 16'h0003;
        rom[159][6] = 16'hFFEE;
        rom[159][7] = 16'h001B;
        rom[159][8] = 16'hFFB9;
        rom[159][9] = 16'h0004;
        rom[159][10] = 16'hFFE8;
        rom[159][11] = 16'h000E;
        rom[159][12] = 16'h0068;
        rom[159][13] = 16'hFFF7;
        rom[159][14] = 16'hFFC2;
        rom[159][15] = 16'h001F;
        rom[159][16] = 16'h000C;
        rom[159][17] = 16'h0020;
        rom[159][18] = 16'h0002;
        rom[159][19] = 16'hFFC8;
        rom[159][20] = 16'hFFEC;
        rom[159][21] = 16'hFFBE;
        rom[159][22] = 16'hFFF5;
        rom[159][23] = 16'hFFF0;
        rom[159][24] = 16'h0010;
        rom[159][25] = 16'hFFA9;
        rom[159][26] = 16'hFFC9;
        rom[159][27] = 16'hFFC1;
        rom[159][28] = 16'h0022;
        rom[159][29] = 16'hFFEE;
        rom[159][30] = 16'hFFCA;
        rom[159][31] = 16'hFFD7;
        rom[159][32] = 16'hFFF6;
        rom[159][33] = 16'hFFF3;
        rom[159][34] = 16'h000F;
        rom[159][35] = 16'hFFDB;
        rom[159][36] = 16'h0018;
        rom[159][37] = 16'h0002;
        rom[159][38] = 16'h0002;
        rom[159][39] = 16'h0005;
        rom[159][40] = 16'h0023;
        rom[159][41] = 16'hFFE6;
        rom[159][42] = 16'hFFB4;
        rom[159][43] = 16'h0002;
        rom[159][44] = 16'h000C;
        rom[159][45] = 16'h0014;
        rom[159][46] = 16'h0012;
        rom[159][47] = 16'hFFDE;
        rom[159][48] = 16'h0034;
        rom[159][49] = 16'hFFFF;
        rom[159][50] = 16'h001D;
        rom[159][51] = 16'hFFC6;
        rom[159][52] = 16'h000B;
        rom[159][53] = 16'h001B;
        rom[159][54] = 16'h0024;
        rom[159][55] = 16'hFFEA;
        rom[159][56] = 16'hFFF6;
        rom[159][57] = 16'hFFEA;
        rom[159][58] = 16'h001F;
        rom[159][59] = 16'hFFD3;
        rom[159][60] = 16'hFFF9;
        rom[159][61] = 16'hFFEE;
        rom[159][62] = 16'hFFF4;
        rom[159][63] = 16'h001F;
        rom[159][64] = 16'h0011;
        rom[159][65] = 16'h0005;
        rom[159][66] = 16'h0004;
        rom[159][67] = 16'hFFCD;
        rom[159][68] = 16'hFFEA;
        rom[159][69] = 16'hFFDE;
        rom[159][70] = 16'hFFE1;
        rom[159][71] = 16'h0002;
        rom[159][72] = 16'hFFC4;
        rom[159][73] = 16'hFFE4;
        rom[159][74] = 16'hFFF3;
        rom[159][75] = 16'hFFED;
        rom[159][76] = 16'h001A;
        rom[159][77] = 16'h002F;
        rom[159][78] = 16'h0015;
        rom[159][79] = 16'h0007;
        rom[159][80] = 16'h0018;
        rom[159][81] = 16'h0013;
        rom[159][82] = 16'hFFFE;
        rom[159][83] = 16'hFFCC;
        rom[159][84] = 16'h000D;
        rom[159][85] = 16'hFFFD;
        rom[159][86] = 16'hFFFB;
        rom[159][87] = 16'h0012;
        rom[159][88] = 16'h000D;
        rom[159][89] = 16'hFFFC;
        rom[159][90] = 16'hFFD5;
        rom[159][91] = 16'h0016;
        rom[159][92] = 16'hFFE5;
        rom[159][93] = 16'h0007;
        rom[159][94] = 16'h002E;
        rom[159][95] = 16'h001A;
        rom[159][96] = 16'h0007;
        rom[159][97] = 16'hFFF3;
        rom[159][98] = 16'hFFBE;
        rom[159][99] = 16'hFFED;
        rom[159][100] = 16'h001C;
        rom[159][101] = 16'h0027;
        rom[159][102] = 16'h0020;
        rom[159][103] = 16'hFFF4;
        rom[159][104] = 16'hFFE1;
        rom[159][105] = 16'hFFF2;
        rom[159][106] = 16'h002E;
        rom[159][107] = 16'h0001;
        rom[159][108] = 16'hFFE8;
        rom[159][109] = 16'h001E;
        rom[159][110] = 16'hFFEE;
        rom[159][111] = 16'hFFEE;
        rom[159][112] = 16'hFFC3;
        rom[159][113] = 16'hFFE1;
        rom[159][114] = 16'hFFCE;
        rom[159][115] = 16'hFFDC;
        rom[159][116] = 16'h001B;
        rom[159][117] = 16'hFFE6;
        rom[159][118] = 16'h002C;
        rom[159][119] = 16'h0002;
        rom[159][120] = 16'h000D;
        rom[159][121] = 16'h001B;
        rom[159][122] = 16'h0003;
        rom[159][123] = 16'h0010;
        rom[159][124] = 16'h0020;
        rom[159][125] = 16'hFFE1;
        rom[159][126] = 16'h0024;
        rom[159][127] = 16'h0002;
        rom[160][0] = 16'hFFED;
        rom[160][1] = 16'h0019;
        rom[160][2] = 16'hFFF8;
        rom[160][3] = 16'h0001;
        rom[160][4] = 16'h0014;
        rom[160][5] = 16'hFFFD;
        rom[160][6] = 16'h000B;
        rom[160][7] = 16'hFFE2;
        rom[160][8] = 16'h000C;
        rom[160][9] = 16'hFFCD;
        rom[160][10] = 16'h0007;
        rom[160][11] = 16'hFFB2;
        rom[160][12] = 16'h0017;
        rom[160][13] = 16'h0021;
        rom[160][14] = 16'h000A;
        rom[160][15] = 16'h0003;
        rom[160][16] = 16'hFFEB;
        rom[160][17] = 16'h001D;
        rom[160][18] = 16'hFFE1;
        rom[160][19] = 16'h000F;
        rom[160][20] = 16'hFFB5;
        rom[160][21] = 16'h0010;
        rom[160][22] = 16'h0024;
        rom[160][23] = 16'hFFDA;
        rom[160][24] = 16'hFFEC;
        rom[160][25] = 16'h000B;
        rom[160][26] = 16'h0006;
        rom[160][27] = 16'h001B;
        rom[160][28] = 16'hFFEA;
        rom[160][29] = 16'hFFFA;
        rom[160][30] = 16'hFFDE;
        rom[160][31] = 16'hFFDA;
        rom[160][32] = 16'h0011;
        rom[160][33] = 16'h0002;
        rom[160][34] = 16'hFFDC;
        rom[160][35] = 16'h0003;
        rom[160][36] = 16'hFFD1;
        rom[160][37] = 16'h000F;
        rom[160][38] = 16'hFFDC;
        rom[160][39] = 16'hFFDC;
        rom[160][40] = 16'h002A;
        rom[160][41] = 16'hFFF6;
        rom[160][42] = 16'hFFFE;
        rom[160][43] = 16'hFFF1;
        rom[160][44] = 16'h000F;
        rom[160][45] = 16'h0029;
        rom[160][46] = 16'hFFB7;
        rom[160][47] = 16'hFFFD;
        rom[160][48] = 16'h0004;
        rom[160][49] = 16'h0014;
        rom[160][50] = 16'h0002;
        rom[160][51] = 16'h0018;
        rom[160][52] = 16'h0016;
        rom[160][53] = 16'h001F;
        rom[160][54] = 16'hFFFF;
        rom[160][55] = 16'h000A;
        rom[160][56] = 16'h000C;
        rom[160][57] = 16'hFFED;
        rom[160][58] = 16'hFFDB;
        rom[160][59] = 16'hFFEC;
        rom[160][60] = 16'h0004;
        rom[160][61] = 16'hFFC9;
        rom[160][62] = 16'h0002;
        rom[160][63] = 16'hFFD7;
        rom[160][64] = 16'hFFF4;
        rom[160][65] = 16'h0015;
        rom[160][66] = 16'h002A;
        rom[160][67] = 16'h0016;
        rom[160][68] = 16'h002E;
        rom[160][69] = 16'hFFF4;
        rom[160][70] = 16'h0016;
        rom[160][71] = 16'h001F;
        rom[160][72] = 16'hFFB8;
        rom[160][73] = 16'h0023;
        rom[160][74] = 16'hFFF8;
        rom[160][75] = 16'hFFE1;
        rom[160][76] = 16'hFFC8;
        rom[160][77] = 16'hFFF4;
        rom[160][78] = 16'h000C;
        rom[160][79] = 16'h0010;
        rom[160][80] = 16'h0004;
        rom[160][81] = 16'hFFDA;
        rom[160][82] = 16'h000C;
        rom[160][83] = 16'hFFEB;
        rom[160][84] = 16'h0014;
        rom[160][85] = 16'hFFD5;
        rom[160][86] = 16'hFFC2;
        rom[160][87] = 16'h0029;
        rom[160][88] = 16'hFFFE;
        rom[160][89] = 16'hFFD7;
        rom[160][90] = 16'hFFF3;
        rom[160][91] = 16'h0019;
        rom[160][92] = 16'h0011;
        rom[160][93] = 16'h0002;
        rom[160][94] = 16'hFFE0;
        rom[160][95] = 16'h0018;
        rom[160][96] = 16'h0015;
        rom[160][97] = 16'h0007;
        rom[160][98] = 16'hFFD0;
        rom[160][99] = 16'hFFE7;
        rom[160][100] = 16'h0009;
        rom[160][101] = 16'hFFE4;
        rom[160][102] = 16'h0000;
        rom[160][103] = 16'h000C;
        rom[160][104] = 16'h002A;
        rom[160][105] = 16'hFFE2;
        rom[160][106] = 16'h0013;
        rom[160][107] = 16'h0013;
        rom[160][108] = 16'hFFF3;
        rom[160][109] = 16'h001A;
        rom[160][110] = 16'h0029;
        rom[160][111] = 16'hFFF4;
        rom[160][112] = 16'hFFC3;
        rom[160][113] = 16'hFFFE;
        rom[160][114] = 16'hFFFE;
        rom[160][115] = 16'h0008;
        rom[160][116] = 16'hFFE5;
        rom[160][117] = 16'hFFF3;
        rom[160][118] = 16'hFFDE;
        rom[160][119] = 16'hFFEE;
        rom[160][120] = 16'h000C;
        rom[160][121] = 16'hFFB8;
        rom[160][122] = 16'hFFD3;
        rom[160][123] = 16'hFFCD;
        rom[160][124] = 16'h0002;
        rom[160][125] = 16'h001A;
        rom[160][126] = 16'h0010;
        rom[160][127] = 16'h0006;
        rom[161][0] = 16'h002E;
        rom[161][1] = 16'hFFA4;
        rom[161][2] = 16'hFFFE;
        rom[161][3] = 16'hFFF5;
        rom[161][4] = 16'hFFFF;
        rom[161][5] = 16'h000A;
        rom[161][6] = 16'hFFE1;
        rom[161][7] = 16'hFFD7;
        rom[161][8] = 16'hFFE1;
        rom[161][9] = 16'hFFDF;
        rom[161][10] = 16'hFFF9;
        rom[161][11] = 16'hFFE9;
        rom[161][12] = 16'hFFFE;
        rom[161][13] = 16'h000A;
        rom[161][14] = 16'hFFE5;
        rom[161][15] = 16'hFFFF;
        rom[161][16] = 16'h0008;
        rom[161][17] = 16'hFFDB;
        rom[161][18] = 16'hFFD8;
        rom[161][19] = 16'hFFB0;
        rom[161][20] = 16'hFFE9;
        rom[161][21] = 16'hFFCA;
        rom[161][22] = 16'hFFFF;
        rom[161][23] = 16'h002A;
        rom[161][24] = 16'h0038;
        rom[161][25] = 16'hFFE5;
        rom[161][26] = 16'hFFB1;
        rom[161][27] = 16'hFFEA;
        rom[161][28] = 16'hFFC5;
        rom[161][29] = 16'hFFBF;
        rom[161][30] = 16'hFFFB;
        rom[161][31] = 16'hFFFF;
        rom[161][32] = 16'hFFF5;
        rom[161][33] = 16'hFFF6;
        rom[161][34] = 16'h0004;
        rom[161][35] = 16'hFFF3;
        rom[161][36] = 16'h0008;
        rom[161][37] = 16'hFFE6;
        rom[161][38] = 16'hFFD2;
        rom[161][39] = 16'hFFD4;
        rom[161][40] = 16'hFFEA;
        rom[161][41] = 16'hFFD8;
        rom[161][42] = 16'hFFCD;
        rom[161][43] = 16'h0026;
        rom[161][44] = 16'hFFE0;
        rom[161][45] = 16'h0015;
        rom[161][46] = 16'hFFD4;
        rom[161][47] = 16'hFFF1;
        rom[161][48] = 16'h001F;
        rom[161][49] = 16'h0016;
        rom[161][50] = 16'h0027;
        rom[161][51] = 16'h001F;
        rom[161][52] = 16'hFFFF;
        rom[161][53] = 16'h0020;
        rom[161][54] = 16'hFFC8;
        rom[161][55] = 16'hFFB8;
        rom[161][56] = 16'hFFE5;
        rom[161][57] = 16'h000A;
        rom[161][58] = 16'hFFEB;
        rom[161][59] = 16'hFFDE;
        rom[161][60] = 16'h0004;
        rom[161][61] = 16'h0017;
        rom[161][62] = 16'hFFC1;
        rom[161][63] = 16'h0009;
        rom[161][64] = 16'hFFF2;
        rom[161][65] = 16'hFFE7;
        rom[161][66] = 16'h0009;
        rom[161][67] = 16'h0021;
        rom[161][68] = 16'h000A;
        rom[161][69] = 16'hFFF2;
        rom[161][70] = 16'h000A;
        rom[161][71] = 16'hFFFC;
        rom[161][72] = 16'h0016;
        rom[161][73] = 16'hFFF9;
        rom[161][74] = 16'h0011;
        rom[161][75] = 16'h0006;
        rom[161][76] = 16'h0028;
        rom[161][77] = 16'hFFEA;
        rom[161][78] = 16'hFFBE;
        rom[161][79] = 16'hFFDA;
        rom[161][80] = 16'hFFDD;
        rom[161][81] = 16'hFFFF;
        rom[161][82] = 16'h0004;
        rom[161][83] = 16'hFFE3;
        rom[161][84] = 16'hFFDC;
        rom[161][85] = 16'h001F;
        rom[161][86] = 16'hFFCC;
        rom[161][87] = 16'h003A;
        rom[161][88] = 16'hFFEA;
        rom[161][89] = 16'hFFF9;
        rom[161][90] = 16'h000C;
        rom[161][91] = 16'h0006;
        rom[161][92] = 16'h0025;
        rom[161][93] = 16'hFFFE;
        rom[161][94] = 16'hFFED;
        rom[161][95] = 16'hFFEF;
        rom[161][96] = 16'hFFED;
        rom[161][97] = 16'h001A;
        rom[161][98] = 16'h0040;
        rom[161][99] = 16'h0028;
        rom[161][100] = 16'h0005;
        rom[161][101] = 16'hFFDC;
        rom[161][102] = 16'h002F;
        rom[161][103] = 16'h000D;
        rom[161][104] = 16'h0001;
        rom[161][105] = 16'h0004;
        rom[161][106] = 16'hFFDC;
        rom[161][107] = 16'h0030;
        rom[161][108] = 16'h0001;
        rom[161][109] = 16'hFFC8;
        rom[161][110] = 16'h0019;
        rom[161][111] = 16'hFFE1;
        rom[161][112] = 16'hFFDC;
        rom[161][113] = 16'hFFEF;
        rom[161][114] = 16'h0013;
        rom[161][115] = 16'hFFA9;
        rom[161][116] = 16'hFFC9;
        rom[161][117] = 16'hFFCF;
        rom[161][118] = 16'h0008;
        rom[161][119] = 16'h000E;
        rom[161][120] = 16'hFFF5;
        rom[161][121] = 16'h0019;
        rom[161][122] = 16'hFFFF;
        rom[161][123] = 16'h0023;
        rom[161][124] = 16'h0013;
        rom[161][125] = 16'h001F;
        rom[161][126] = 16'h0000;
        rom[161][127] = 16'hFFF1;
        rom[162][0] = 16'hFFC1;
        rom[162][1] = 16'hFFF7;
        rom[162][2] = 16'h0004;
        rom[162][3] = 16'h002B;
        rom[162][4] = 16'hFFC5;
        rom[162][5] = 16'hFFBA;
        rom[162][6] = 16'hFFE3;
        rom[162][7] = 16'hFFDE;
        rom[162][8] = 16'h0002;
        rom[162][9] = 16'hFFEA;
        rom[162][10] = 16'h000C;
        rom[162][11] = 16'hFFFB;
        rom[162][12] = 16'hFFE8;
        rom[162][13] = 16'h0028;
        rom[162][14] = 16'hFFF5;
        rom[162][15] = 16'h000D;
        rom[162][16] = 16'hFFFE;
        rom[162][17] = 16'h0012;
        rom[162][18] = 16'h0017;
        rom[162][19] = 16'h0024;
        rom[162][20] = 16'h0011;
        rom[162][21] = 16'h001D;
        rom[162][22] = 16'hFFF4;
        rom[162][23] = 16'hFFF8;
        rom[162][24] = 16'hFFE2;
        rom[162][25] = 16'h003B;
        rom[162][26] = 16'h0001;
        rom[162][27] = 16'h002A;
        rom[162][28] = 16'h000B;
        rom[162][29] = 16'h0033;
        rom[162][30] = 16'hFFD5;
        rom[162][31] = 16'h001F;
        rom[162][32] = 16'h000D;
        rom[162][33] = 16'hFFEC;
        rom[162][34] = 16'hFFEA;
        rom[162][35] = 16'hFFF4;
        rom[162][36] = 16'hFFE9;
        rom[162][37] = 16'h0010;
        rom[162][38] = 16'hFFE7;
        rom[162][39] = 16'hFFDF;
        rom[162][40] = 16'hFFE3;
        rom[162][41] = 16'hFFD2;
        rom[162][42] = 16'hFFDB;
        rom[162][43] = 16'h0024;
        rom[162][44] = 16'hFFDB;
        rom[162][45] = 16'h0016;
        rom[162][46] = 16'hFFE0;
        rom[162][47] = 16'h0002;
        rom[162][48] = 16'hFFCA;
        rom[162][49] = 16'hFFE0;
        rom[162][50] = 16'hFFFE;
        rom[162][51] = 16'hFFE4;
        rom[162][52] = 16'hFFEF;
        rom[162][53] = 16'h002A;
        rom[162][54] = 16'h0002;
        rom[162][55] = 16'hFFE8;
        rom[162][56] = 16'hFFF1;
        rom[162][57] = 16'hFFEF;
        rom[162][58] = 16'hFFE4;
        rom[162][59] = 16'h0029;
        rom[162][60] = 16'h0002;
        rom[162][61] = 16'h0007;
        rom[162][62] = 16'hFFDE;
        rom[162][63] = 16'hFFDD;
        rom[162][64] = 16'h0003;
        rom[162][65] = 16'hFFCB;
        rom[162][66] = 16'hFFFC;
        rom[162][67] = 16'hFFF2;
        rom[162][68] = 16'hFFE5;
        rom[162][69] = 16'hFFFA;
        rom[162][70] = 16'h000A;
        rom[162][71] = 16'h0011;
        rom[162][72] = 16'hFFFE;
        rom[162][73] = 16'hFFD2;
        rom[162][74] = 16'hFFD1;
        rom[162][75] = 16'hFFDC;
        rom[162][76] = 16'hFFEF;
        rom[162][77] = 16'hFFC3;
        rom[162][78] = 16'h0017;
        rom[162][79] = 16'hFFC9;
        rom[162][80] = 16'h001F;
        rom[162][81] = 16'hFFF5;
        rom[162][82] = 16'h0015;
        rom[162][83] = 16'hFFFF;
        rom[162][84] = 16'hFFCE;
        rom[162][85] = 16'hFFF0;
        rom[162][86] = 16'hFFD7;
        rom[162][87] = 16'hFFEF;
        rom[162][88] = 16'h0012;
        rom[162][89] = 16'hFFFA;
        rom[162][90] = 16'h001E;
        rom[162][91] = 16'h001B;
        rom[162][92] = 16'hFFDF;
        rom[162][93] = 16'hFFF4;
        rom[162][94] = 16'hFFEB;
        rom[162][95] = 16'hFFC8;
        rom[162][96] = 16'hFFD9;
        rom[162][97] = 16'hFFDB;
        rom[162][98] = 16'hFFF7;
        rom[162][99] = 16'hFFE6;
        rom[162][100] = 16'hFFD7;
        rom[162][101] = 16'hFFD0;
        rom[162][102] = 16'h0005;
        rom[162][103] = 16'hFFF8;
        rom[162][104] = 16'h0011;
        rom[162][105] = 16'hFFF9;
        rom[162][106] = 16'hFFF2;
        rom[162][107] = 16'hFFE1;
        rom[162][108] = 16'hFFCA;
        rom[162][109] = 16'h0007;
        rom[162][110] = 16'hFFED;
        rom[162][111] = 16'h0006;
        rom[162][112] = 16'hFFFC;
        rom[162][113] = 16'h001C;
        rom[162][114] = 16'hFFFA;
        rom[162][115] = 16'h0000;
        rom[162][116] = 16'hFFDD;
        rom[162][117] = 16'h0003;
        rom[162][118] = 16'hFFE4;
        rom[162][119] = 16'hFFDA;
        rom[162][120] = 16'hFFF2;
        rom[162][121] = 16'hFFF2;
        rom[162][122] = 16'hFFF4;
        rom[162][123] = 16'hFFEF;
        rom[162][124] = 16'h001C;
        rom[162][125] = 16'hFFD4;
        rom[162][126] = 16'h0012;
        rom[162][127] = 16'hFFDD;
        rom[163][0] = 16'hFFC0;
        rom[163][1] = 16'h000C;
        rom[163][2] = 16'hFFE5;
        rom[163][3] = 16'h0002;
        rom[163][4] = 16'h0013;
        rom[163][5] = 16'h0015;
        rom[163][6] = 16'hFFFD;
        rom[163][7] = 16'h0016;
        rom[163][8] = 16'h0016;
        rom[163][9] = 16'hFFE4;
        rom[163][10] = 16'h0000;
        rom[163][11] = 16'hFFE5;
        rom[163][12] = 16'h0007;
        rom[163][13] = 16'hFFD5;
        rom[163][14] = 16'h0004;
        rom[163][15] = 16'h0008;
        rom[163][16] = 16'h0017;
        rom[163][17] = 16'h0002;
        rom[163][18] = 16'hFFC5;
        rom[163][19] = 16'hFFF4;
        rom[163][20] = 16'hFFE7;
        rom[163][21] = 16'hFFF8;
        rom[163][22] = 16'hFFCD;
        rom[163][23] = 16'h0017;
        rom[163][24] = 16'hFFE3;
        rom[163][25] = 16'hFFD2;
        rom[163][26] = 16'hFFEE;
        rom[163][27] = 16'h0005;
        rom[163][28] = 16'hFFFD;
        rom[163][29] = 16'hFFFD;
        rom[163][30] = 16'h002E;
        rom[163][31] = 16'h000B;
        rom[163][32] = 16'hFFFE;
        rom[163][33] = 16'hFFC6;
        rom[163][34] = 16'hFFFC;
        rom[163][35] = 16'hFFFE;
        rom[163][36] = 16'h0016;
        rom[163][37] = 16'hFFC5;
        rom[163][38] = 16'hFFD8;
        rom[163][39] = 16'hFFF1;
        rom[163][40] = 16'h0031;
        rom[163][41] = 16'hFFDB;
        rom[163][42] = 16'hFFE4;
        rom[163][43] = 16'hFFED;
        rom[163][44] = 16'h0002;
        rom[163][45] = 16'hFFE1;
        rom[163][46] = 16'h0000;
        rom[163][47] = 16'hFFEF;
        rom[163][48] = 16'hFFED;
        rom[163][49] = 16'h0028;
        rom[163][50] = 16'hFFE1;
        rom[163][51] = 16'hFFF9;
        rom[163][52] = 16'h0019;
        rom[163][53] = 16'h0024;
        rom[163][54] = 16'h0002;
        rom[163][55] = 16'h001F;
        rom[163][56] = 16'h001E;
        rom[163][57] = 16'h0012;
        rom[163][58] = 16'hFFF5;
        rom[163][59] = 16'h000D;
        rom[163][60] = 16'h0025;
        rom[163][61] = 16'h0028;
        rom[163][62] = 16'hFFB0;
        rom[163][63] = 16'h0000;
        rom[163][64] = 16'h0002;
        rom[163][65] = 16'hFFE9;
        rom[163][66] = 16'h002E;
        rom[163][67] = 16'h0011;
        rom[163][68] = 16'h0002;
        rom[163][69] = 16'h001F;
        rom[163][70] = 16'h0013;
        rom[163][71] = 16'hFFE5;
        rom[163][72] = 16'hFFE5;
        rom[163][73] = 16'h0010;
        rom[163][74] = 16'hFFF1;
        rom[163][75] = 16'hFFDF;
        rom[163][76] = 16'hFFDC;
        rom[163][77] = 16'h0018;
        rom[163][78] = 16'hFFD2;
        rom[163][79] = 16'h0022;
        rom[163][80] = 16'hFFEE;
        rom[163][81] = 16'hFFC2;
        rom[163][82] = 16'h0027;
        rom[163][83] = 16'h000B;
        rom[163][84] = 16'hFFEF;
        rom[163][85] = 16'h000F;
        rom[163][86] = 16'h0018;
        rom[163][87] = 16'h000F;
        rom[163][88] = 16'hFFCD;
        rom[163][89] = 16'hFFF9;
        rom[163][90] = 16'h0038;
        rom[163][91] = 16'hFFDE;
        rom[163][92] = 16'hFFE1;
        rom[163][93] = 16'h0014;
        rom[163][94] = 16'hFFEA;
        rom[163][95] = 16'hFFE6;
        rom[163][96] = 16'h0006;
        rom[163][97] = 16'hFFEB;
        rom[163][98] = 16'h0005;
        rom[163][99] = 16'h000C;
        rom[163][100] = 16'hFFF8;
        rom[163][101] = 16'hFFBC;
        rom[163][102] = 16'hFFE1;
        rom[163][103] = 16'hFFCD;
        rom[163][104] = 16'h0017;
        rom[163][105] = 16'h0015;
        rom[163][106] = 16'h000F;
        rom[163][107] = 16'hFFF0;
        rom[163][108] = 16'hFFF4;
        rom[163][109] = 16'hFFF8;
        rom[163][110] = 16'h001D;
        rom[163][111] = 16'h0002;
        rom[163][112] = 16'hFFD0;
        rom[163][113] = 16'h001A;
        rom[163][114] = 16'h000D;
        rom[163][115] = 16'h0029;
        rom[163][116] = 16'hFFEF;
        rom[163][117] = 16'h0003;
        rom[163][118] = 16'hFFFC;
        rom[163][119] = 16'hFFA2;
        rom[163][120] = 16'h0002;
        rom[163][121] = 16'h002E;
        rom[163][122] = 16'h0002;
        rom[163][123] = 16'hFFF2;
        rom[163][124] = 16'hFFFA;
        rom[163][125] = 16'h0008;
        rom[163][126] = 16'h0018;
        rom[163][127] = 16'hFFFA;
        rom[164][0] = 16'h0002;
        rom[164][1] = 16'h0002;
        rom[164][2] = 16'h0010;
        rom[164][3] = 16'h0007;
        rom[164][4] = 16'h0028;
        rom[164][5] = 16'h0006;
        rom[164][6] = 16'hFFE3;
        rom[164][7] = 16'hFFF4;
        rom[164][8] = 16'h0023;
        rom[164][9] = 16'hFFE5;
        rom[164][10] = 16'h003B;
        rom[164][11] = 16'h0029;
        rom[164][12] = 16'h0006;
        rom[164][13] = 16'h0017;
        rom[164][14] = 16'h0024;
        rom[164][15] = 16'hFFF7;
        rom[164][16] = 16'h0007;
        rom[164][17] = 16'hFFD2;
        rom[164][18] = 16'hFFF6;
        rom[164][19] = 16'hFFEF;
        rom[164][20] = 16'h0007;
        rom[164][21] = 16'hFFE7;
        rom[164][22] = 16'hFFE4;
        rom[164][23] = 16'h0024;
        rom[164][24] = 16'hFFB5;
        rom[164][25] = 16'h0005;
        rom[164][26] = 16'h0000;
        rom[164][27] = 16'h0015;
        rom[164][28] = 16'h0015;
        rom[164][29] = 16'hFFE5;
        rom[164][30] = 16'h0027;
        rom[164][31] = 16'hFFE9;
        rom[164][32] = 16'h0007;
        rom[164][33] = 16'hFFCE;
        rom[164][34] = 16'h001E;
        rom[164][35] = 16'hFFDB;
        rom[164][36] = 16'hFFEA;
        rom[164][37] = 16'hFFD7;
        rom[164][38] = 16'hFFA7;
        rom[164][39] = 16'hFFE7;
        rom[164][40] = 16'h0034;
        rom[164][41] = 16'hFFFD;
        rom[164][42] = 16'h0016;
        rom[164][43] = 16'h000C;
        rom[164][44] = 16'hFFE3;
        rom[164][45] = 16'hFFE2;
        rom[164][46] = 16'hFFFF;
        rom[164][47] = 16'hFFFB;
        rom[164][48] = 16'h000D;
        rom[164][49] = 16'h000C;
        rom[164][50] = 16'hFFEF;
        rom[164][51] = 16'h0018;
        rom[164][52] = 16'h0000;
        rom[164][53] = 16'h0029;
        rom[164][54] = 16'h0002;
        rom[164][55] = 16'hFFF6;
        rom[164][56] = 16'hFFF3;
        rom[164][57] = 16'hFFF9;
        rom[164][58] = 16'hFFCD;
        rom[164][59] = 16'h001B;
        rom[164][60] = 16'h0009;
        rom[164][61] = 16'hFFCA;
        rom[164][62] = 16'h0017;
        rom[164][63] = 16'hFFD2;
        rom[164][64] = 16'hFFE5;
        rom[164][65] = 16'h000D;
        rom[164][66] = 16'h0025;
        rom[164][67] = 16'h0023;
        rom[164][68] = 16'hFFDC;
        rom[164][69] = 16'h001B;
        rom[164][70] = 16'hFFD2;
        rom[164][71] = 16'h000B;
        rom[164][72] = 16'h0015;
        rom[164][73] = 16'h0025;
        rom[164][74] = 16'hFFDA;
        rom[164][75] = 16'hFFBA;
        rom[164][76] = 16'hFFD7;
        rom[164][77] = 16'hFFFA;
        rom[164][78] = 16'h0003;
        rom[164][79] = 16'hFFFD;
        rom[164][80] = 16'hFFE3;
        rom[164][81] = 16'hFFAC;
        rom[164][82] = 16'h0013;
        rom[164][83] = 16'hFFCD;
        rom[164][84] = 16'hFFC4;
        rom[164][85] = 16'h0008;
        rom[164][86] = 16'h000B;
        rom[164][87] = 16'h0028;
        rom[164][88] = 16'hFFB7;
        rom[164][89] = 16'h000F;
        rom[164][90] = 16'h0006;
        rom[164][91] = 16'h0041;
        rom[164][92] = 16'h000C;
        rom[164][93] = 16'hFFD7;
        rom[164][94] = 16'h0005;
        rom[164][95] = 16'hFFD7;
        rom[164][96] = 16'h0001;
        rom[164][97] = 16'h0020;
        rom[164][98] = 16'h001F;
        rom[164][99] = 16'hFFE6;
        rom[164][100] = 16'h0025;
        rom[164][101] = 16'hFFD5;
        rom[164][102] = 16'hFFF4;
        rom[164][103] = 16'hFFCC;
        rom[164][104] = 16'h0009;
        rom[164][105] = 16'hFFC1;
        rom[164][106] = 16'hFFCA;
        rom[164][107] = 16'hFFF4;
        rom[164][108] = 16'h0041;
        rom[164][109] = 16'hFFD5;
        rom[164][110] = 16'h0014;
        rom[164][111] = 16'h0005;
        rom[164][112] = 16'hFFEA;
        rom[164][113] = 16'hFFF9;
        rom[164][114] = 16'hFFF4;
        rom[164][115] = 16'hFFFF;
        rom[164][116] = 16'hFFF4;
        rom[164][117] = 16'h0016;
        rom[164][118] = 16'hFFE2;
        rom[164][119] = 16'hFFBF;
        rom[164][120] = 16'h000C;
        rom[164][121] = 16'h001C;
        rom[164][122] = 16'h0016;
        rom[164][123] = 16'h000D;
        rom[164][124] = 16'h0023;
        rom[164][125] = 16'h001A;
        rom[164][126] = 16'h0014;
        rom[164][127] = 16'h0014;
        rom[165][0] = 16'h000C;
        rom[165][1] = 16'h0018;
        rom[165][2] = 16'hFFE5;
        rom[165][3] = 16'h0016;
        rom[165][4] = 16'h0002;
        rom[165][5] = 16'hFFE0;
        rom[165][6] = 16'hFFF7;
        rom[165][7] = 16'h0011;
        rom[165][8] = 16'hFFF4;
        rom[165][9] = 16'h0016;
        rom[165][10] = 16'h002B;
        rom[165][11] = 16'hFFF1;
        rom[165][12] = 16'h002A;
        rom[165][13] = 16'h0007;
        rom[165][14] = 16'h0013;
        rom[165][15] = 16'hFFFE;
        rom[165][16] = 16'h0021;
        rom[165][17] = 16'hFFF7;
        rom[165][18] = 16'hFFF6;
        rom[165][19] = 16'hFFE6;
        rom[165][20] = 16'hFFD6;
        rom[165][21] = 16'h000C;
        rom[165][22] = 16'h0028;
        rom[165][23] = 16'h0011;
        rom[165][24] = 16'hFFF4;
        rom[165][25] = 16'hFFD2;
        rom[165][26] = 16'hFFFD;
        rom[165][27] = 16'hFFBF;
        rom[165][28] = 16'h0024;
        rom[165][29] = 16'hFFFC;
        rom[165][30] = 16'hFFF4;
        rom[165][31] = 16'h0012;
        rom[165][32] = 16'hFFF5;
        rom[165][33] = 16'hFFF3;
        rom[165][34] = 16'h0023;
        rom[165][35] = 16'h0005;
        rom[165][36] = 16'h0019;
        rom[165][37] = 16'hFFE6;
        rom[165][38] = 16'h000C;
        rom[165][39] = 16'h0004;
        rom[165][40] = 16'hFFF0;
        rom[165][41] = 16'hFFE5;
        rom[165][42] = 16'h0021;
        rom[165][43] = 16'h0023;
        rom[165][44] = 16'h0047;
        rom[165][45] = 16'hFFD5;
        rom[165][46] = 16'h001C;
        rom[165][47] = 16'h000B;
        rom[165][48] = 16'hFFF6;
        rom[165][49] = 16'hFFE1;
        rom[165][50] = 16'h0008;
        rom[165][51] = 16'h001B;
        rom[165][52] = 16'h0033;
        rom[165][53] = 16'hFFCF;
        rom[165][54] = 16'hFFD8;
        rom[165][55] = 16'hFFC4;
        rom[165][56] = 16'hFFC1;
        rom[165][57] = 16'hFFF4;
        rom[165][58] = 16'h0017;
        rom[165][59] = 16'hFFD5;
        rom[165][60] = 16'h0019;
        rom[165][61] = 16'h001E;
        rom[165][62] = 16'hFFC3;
        rom[165][63] = 16'hFFDC;
        rom[165][64] = 16'h0029;
        rom[165][65] = 16'h0016;
        rom[165][66] = 16'hFFF5;
        rom[165][67] = 16'hFFF1;
        rom[165][68] = 16'hFFEF;
        rom[165][69] = 16'h001F;
        rom[165][70] = 16'h0002;
        rom[165][71] = 16'hFFEA;
        rom[165][72] = 16'hFFF0;
        rom[165][73] = 16'hFFEB;
        rom[165][74] = 16'h000E;
        rom[165][75] = 16'hFFE7;
        rom[165][76] = 16'hFFDC;
        rom[165][77] = 16'hFFEC;
        rom[165][78] = 16'hFFE9;
        rom[165][79] = 16'hFFFE;
        rom[165][80] = 16'hFFE5;
        rom[165][81] = 16'h0013;
        rom[165][82] = 16'hFFE3;
        rom[165][83] = 16'hFFF0;
        rom[165][84] = 16'h0007;
        rom[165][85] = 16'hFFE5;
        rom[165][86] = 16'hFFFF;
        rom[165][87] = 16'h0002;
        rom[165][88] = 16'hFFE6;
        rom[165][89] = 16'hFFB6;
        rom[165][90] = 16'hFFF5;
        rom[165][91] = 16'h003A;
        rom[165][92] = 16'h0009;
        rom[165][93] = 16'hFFEC;
        rom[165][94] = 16'h0016;
        rom[165][95] = 16'hFFE4;
        rom[165][96] = 16'hFFE0;
        rom[165][97] = 16'hFFAB;
        rom[165][98] = 16'h000A;
        rom[165][99] = 16'h0033;
        rom[165][100] = 16'hFFD5;
        rom[165][101] = 16'h0019;
        rom[165][102] = 16'h0007;
        rom[165][103] = 16'hFFFC;
        rom[165][104] = 16'h001D;
        rom[165][105] = 16'hFFF4;
        rom[165][106] = 16'h0032;
        rom[165][107] = 16'hFFFD;
        rom[165][108] = 16'h0000;
        rom[165][109] = 16'h000D;
        rom[165][110] = 16'hFFFC;
        rom[165][111] = 16'h000C;
        rom[165][112] = 16'hFFCF;
        rom[165][113] = 16'hFFEB;
        rom[165][114] = 16'h0024;
        rom[165][115] = 16'h0007;
        rom[165][116] = 16'h0018;
        rom[165][117] = 16'h0002;
        rom[165][118] = 16'hFFEA;
        rom[165][119] = 16'h0000;
        rom[165][120] = 16'h0018;
        rom[165][121] = 16'hFFD1;
        rom[165][122] = 16'hFFE1;
        rom[165][123] = 16'h003F;
        rom[165][124] = 16'h0009;
        rom[165][125] = 16'h001F;
        rom[165][126] = 16'h000A;
        rom[165][127] = 16'h0001;
        rom[166][0] = 16'hFFE6;
        rom[166][1] = 16'h001D;
        rom[166][2] = 16'h0008;
        rom[166][3] = 16'hFFDB;
        rom[166][4] = 16'hFFDE;
        rom[166][5] = 16'hFFF4;
        rom[166][6] = 16'h0005;
        rom[166][7] = 16'h0008;
        rom[166][8] = 16'h000C;
        rom[166][9] = 16'hFFED;
        rom[166][10] = 16'hFFC9;
        rom[166][11] = 16'hFFC8;
        rom[166][12] = 16'h0008;
        rom[166][13] = 16'hFFF1;
        rom[166][14] = 16'hFFEF;
        rom[166][15] = 16'hFFE9;
        rom[166][16] = 16'h0000;
        rom[166][17] = 16'hFFFE;
        rom[166][18] = 16'h000C;
        rom[166][19] = 16'hFFF8;
        rom[166][20] = 16'h000C;
        rom[166][21] = 16'hFFDB;
        rom[166][22] = 16'h0002;
        rom[166][23] = 16'hFFA6;
        rom[166][24] = 16'hFFFE;
        rom[166][25] = 16'h0029;
        rom[166][26] = 16'h001B;
        rom[166][27] = 16'hFFD5;
        rom[166][28] = 16'hFFA9;
        rom[166][29] = 16'hFFE5;
        rom[166][30] = 16'h0002;
        rom[166][31] = 16'h0007;
        rom[166][32] = 16'hFFF9;
        rom[166][33] = 16'hFFF2;
        rom[166][34] = 16'hFFC6;
        rom[166][35] = 16'hFFD1;
        rom[166][36] = 16'h0027;
        rom[166][37] = 16'h0005;
        rom[166][38] = 16'h000F;
        rom[166][39] = 16'hFFCA;
        rom[166][40] = 16'hFFEC;
        rom[166][41] = 16'hFFFC;
        rom[166][42] = 16'hFFD2;
        rom[166][43] = 16'h001F;
        rom[166][44] = 16'hFFB9;
        rom[166][45] = 16'hFFED;
        rom[166][46] = 16'h0025;
        rom[166][47] = 16'h0036;
        rom[166][48] = 16'h0008;
        rom[166][49] = 16'h0029;
        rom[166][50] = 16'hFFF4;
        rom[166][51] = 16'hFFF1;
        rom[166][52] = 16'hFFFF;
        rom[166][53] = 16'h0002;
        rom[166][54] = 16'h000C;
        rom[166][55] = 16'h0003;
        rom[166][56] = 16'hFFFF;
        rom[166][57] = 16'hFFEC;
        rom[166][58] = 16'h002E;
        rom[166][59] = 16'h0008;
        rom[166][60] = 16'hFFC1;
        rom[166][61] = 16'hFFCE;
        rom[166][62] = 16'h0020;
        rom[166][63] = 16'h001E;
        rom[166][64] = 16'h0003;
        rom[166][65] = 16'h000C;
        rom[166][66] = 16'hFFFC;
        rom[166][67] = 16'hFFF4;
        rom[166][68] = 16'h001D;
        rom[166][69] = 16'h0009;
        rom[166][70] = 16'h000B;
        rom[166][71] = 16'h000F;
        rom[166][72] = 16'hFFFA;
        rom[166][73] = 16'hFFE9;
        rom[166][74] = 16'hFFFB;
        rom[166][75] = 16'h0026;
        rom[166][76] = 16'hFFF8;
        rom[166][77] = 16'h0017;
        rom[166][78] = 16'hFFD1;
        rom[166][79] = 16'h0014;
        rom[166][80] = 16'h003C;
        rom[166][81] = 16'h0012;
        rom[166][82] = 16'h0007;
        rom[166][83] = 16'hFFF9;
        rom[166][84] = 16'hFFF5;
        rom[166][85] = 16'h0000;
        rom[166][86] = 16'hFFF5;
        rom[166][87] = 16'h0002;
        rom[166][88] = 16'h0012;
        rom[166][89] = 16'hFFF4;
        rom[166][90] = 16'h001F;
        rom[166][91] = 16'h0032;
        rom[166][92] = 16'h0004;
        rom[166][93] = 16'hFFB5;
        rom[166][94] = 16'h001E;
        rom[166][95] = 16'hFFE0;
        rom[166][96] = 16'hFFFE;
        rom[166][97] = 16'h002F;
        rom[166][98] = 16'hFFF4;
        rom[166][99] = 16'hFFF1;
        rom[166][100] = 16'h0061;
        rom[166][101] = 16'hFFE3;
        rom[166][102] = 16'h0011;
        rom[166][103] = 16'h0003;
        rom[166][104] = 16'hFFE2;
        rom[166][105] = 16'h000B;
        rom[166][106] = 16'h0000;
        rom[166][107] = 16'hFFDC;
        rom[166][108] = 16'hFFEA;
        rom[166][109] = 16'hFFE4;
        rom[166][110] = 16'hFFE8;
        rom[166][111] = 16'hFFE9;
        rom[166][112] = 16'hFFE4;
        rom[166][113] = 16'h0036;
        rom[166][114] = 16'hFFEF;
        rom[166][115] = 16'hFFA9;
        rom[166][116] = 16'h0009;
        rom[166][117] = 16'hFFD0;
        rom[166][118] = 16'h001B;
        rom[166][119] = 16'hFFFA;
        rom[166][120] = 16'hFFB8;
        rom[166][121] = 16'hFFE3;
        rom[166][122] = 16'hFFE7;
        rom[166][123] = 16'h001C;
        rom[166][124] = 16'h0008;
        rom[166][125] = 16'hFFEF;
        rom[166][126] = 16'h0001;
        rom[166][127] = 16'hFFFF;
        rom[167][0] = 16'hFFE9;
        rom[167][1] = 16'h0006;
        rom[167][2] = 16'hFFF3;
        rom[167][3] = 16'hFFFD;
        rom[167][4] = 16'hFFED;
        rom[167][5] = 16'hFFFB;
        rom[167][6] = 16'hFFFB;
        rom[167][7] = 16'hFFFF;
        rom[167][8] = 16'hFFEF;
        rom[167][9] = 16'h000C;
        rom[167][10] = 16'h0009;
        rom[167][11] = 16'h0000;
        rom[167][12] = 16'h0004;
        rom[167][13] = 16'hFFF3;
        rom[167][14] = 16'h0018;
        rom[167][15] = 16'h0006;
        rom[167][16] = 16'hFFF3;
        rom[167][17] = 16'hFFF2;
        rom[167][18] = 16'hFFE7;
        rom[167][19] = 16'hFFCE;
        rom[167][20] = 16'hFFE5;
        rom[167][21] = 16'hFFF2;
        rom[167][22] = 16'hFFDD;
        rom[167][23] = 16'hFFFC;
        rom[167][24] = 16'h0005;
        rom[167][25] = 16'hFFDE;
        rom[167][26] = 16'hFFF1;
        rom[167][27] = 16'hFFAD;
        rom[167][28] = 16'hFFFE;
        rom[167][29] = 16'hFFFB;
        rom[167][30] = 16'hFFD6;
        rom[167][31] = 16'hFFEF;
        rom[167][32] = 16'hFFE1;
        rom[167][33] = 16'h0008;
        rom[167][34] = 16'hFFDE;
        rom[167][35] = 16'h001F;
        rom[167][36] = 16'hFFFB;
        rom[167][37] = 16'hFFF7;
        rom[167][38] = 16'hFFF9;
        rom[167][39] = 16'hFFF7;
        rom[167][40] = 16'hFFFA;
        rom[167][41] = 16'h001C;
        rom[167][42] = 16'h0006;
        rom[167][43] = 16'h001F;
        rom[167][44] = 16'hFFE8;
        rom[167][45] = 16'h0021;
        rom[167][46] = 16'h0003;
        rom[167][47] = 16'h0027;
        rom[167][48] = 16'h001A;
        rom[167][49] = 16'hFFFA;
        rom[167][50] = 16'hFFFF;
        rom[167][51] = 16'hFFBE;
        rom[167][52] = 16'hFFF5;
        rom[167][53] = 16'h0016;
        rom[167][54] = 16'hFFFB;
        rom[167][55] = 16'hFFCC;
        rom[167][56] = 16'h0007;
        rom[167][57] = 16'hFFE5;
        rom[167][58] = 16'hFFFE;
        rom[167][59] = 16'hFFE9;
        rom[167][60] = 16'h000E;
        rom[167][61] = 16'hFFE9;
        rom[167][62] = 16'h0019;
        rom[167][63] = 16'hFFF6;
        rom[167][64] = 16'h0007;
        rom[167][65] = 16'h000C;
        rom[167][66] = 16'hFFF4;
        rom[167][67] = 16'hFFF2;
        rom[167][68] = 16'hFFF3;
        rom[167][69] = 16'hFFDE;
        rom[167][70] = 16'hFFED;
        rom[167][71] = 16'h000F;
        rom[167][72] = 16'h0005;
        rom[167][73] = 16'hFFD2;
        rom[167][74] = 16'h0002;
        rom[167][75] = 16'hFFFF;
        rom[167][76] = 16'h000A;
        rom[167][77] = 16'h0030;
        rom[167][78] = 16'hFFBF;
        rom[167][79] = 16'h0004;
        rom[167][80] = 16'h0007;
        rom[167][81] = 16'h0014;
        rom[167][82] = 16'hFFD7;
        rom[167][83] = 16'hFFF7;
        rom[167][84] = 16'hFFFA;
        rom[167][85] = 16'hFFF8;
        rom[167][86] = 16'h001D;
        rom[167][87] = 16'hFFE3;
        rom[167][88] = 16'hFFBA;
        rom[167][89] = 16'hFFE4;
        rom[167][90] = 16'hFFC3;
        rom[167][91] = 16'hFFD6;
        rom[167][92] = 16'hFFE7;
        rom[167][93] = 16'hFFD9;
        rom[167][94] = 16'h0011;
        rom[167][95] = 16'hFFCC;
        rom[167][96] = 16'hFFEC;
        rom[167][97] = 16'h002D;
        rom[167][98] = 16'hFFF5;
        rom[167][99] = 16'hFFE1;
        rom[167][100] = 16'hFFE2;
        rom[167][101] = 16'h0009;
        rom[167][102] = 16'h0034;
        rom[167][103] = 16'h0016;
        rom[167][104] = 16'hFFD2;
        rom[167][105] = 16'hFFC2;
        rom[167][106] = 16'hFFF2;
        rom[167][107] = 16'h0010;
        rom[167][108] = 16'hFFC9;
        rom[167][109] = 16'h002E;
        rom[167][110] = 16'h0005;
        rom[167][111] = 16'hFFC7;
        rom[167][112] = 16'hFFD7;
        rom[167][113] = 16'hFFD3;
        rom[167][114] = 16'h0013;
        rom[167][115] = 16'hFFDE;
        rom[167][116] = 16'hFFFA;
        rom[167][117] = 16'h001F;
        rom[167][118] = 16'hFFFD;
        rom[167][119] = 16'h001A;
        rom[167][120] = 16'h0002;
        rom[167][121] = 16'hFFE3;
        rom[167][122] = 16'h000A;
        rom[167][123] = 16'hFFF6;
        rom[167][124] = 16'hFFF4;
        rom[167][125] = 16'hFFE5;
        rom[167][126] = 16'hFFEA;
        rom[167][127] = 16'hFFCB;
        rom[168][0] = 16'h000F;
        rom[168][1] = 16'h0014;
        rom[168][2] = 16'hFFFA;
        rom[168][3] = 16'hFFBE;
        rom[168][4] = 16'hFFF9;
        rom[168][5] = 16'h0001;
        rom[168][6] = 16'h0030;
        rom[168][7] = 16'hFFD9;
        rom[168][8] = 16'hFFC9;
        rom[168][9] = 16'hFFE2;
        rom[168][10] = 16'hFFF3;
        rom[168][11] = 16'h0025;
        rom[168][12] = 16'hFFF0;
        rom[168][13] = 16'hFFE9;
        rom[168][14] = 16'h0004;
        rom[168][15] = 16'hFFD5;
        rom[168][16] = 16'h0022;
        rom[168][17] = 16'hFFD9;
        rom[168][18] = 16'hFFEF;
        rom[168][19] = 16'hFFD2;
        rom[168][20] = 16'h001B;
        rom[168][21] = 16'hFFFB;
        rom[168][22] = 16'h002C;
        rom[168][23] = 16'h0016;
        rom[168][24] = 16'h001B;
        rom[168][25] = 16'hFFFA;
        rom[168][26] = 16'h0015;
        rom[168][27] = 16'h0017;
        rom[168][28] = 16'hFFEA;
        rom[168][29] = 16'hFFE0;
        rom[168][30] = 16'h000C;
        rom[168][31] = 16'hFFE2;
        rom[168][32] = 16'hFFD2;
        rom[168][33] = 16'h0010;
        rom[168][34] = 16'hFFFF;
        rom[168][35] = 16'hFFE6;
        rom[168][36] = 16'h0026;
        rom[168][37] = 16'h0008;
        rom[168][38] = 16'h0002;
        rom[168][39] = 16'hFFD0;
        rom[168][40] = 16'h0009;
        rom[168][41] = 16'h0003;
        rom[168][42] = 16'hFFEA;
        rom[168][43] = 16'h0006;
        rom[168][44] = 16'hFFBB;
        rom[168][45] = 16'hFFC1;
        rom[168][46] = 16'hFFFF;
        rom[168][47] = 16'h0008;
        rom[168][48] = 16'h0011;
        rom[168][49] = 16'h0004;
        rom[168][50] = 16'h0012;
        rom[168][51] = 16'h0002;
        rom[168][52] = 16'h0002;
        rom[168][53] = 16'hFFEF;
        rom[168][54] = 16'hFFE3;
        rom[168][55] = 16'hFFF4;
        rom[168][56] = 16'h000C;
        rom[168][57] = 16'h0020;
        rom[168][58] = 16'h0019;
        rom[168][59] = 16'hFFFD;
        rom[168][60] = 16'h0000;
        rom[168][61] = 16'hFFE6;
        rom[168][62] = 16'h001A;
        rom[168][63] = 16'hFFEE;
        rom[168][64] = 16'hFFFE;
        rom[168][65] = 16'hFFE3;
        rom[168][66] = 16'hFFDC;
        rom[168][67] = 16'h0013;
        rom[168][68] = 16'hFFF0;
        rom[168][69] = 16'hFFE8;
        rom[168][70] = 16'hFFF4;
        rom[168][71] = 16'h0021;
        rom[168][72] = 16'h000F;
        rom[168][73] = 16'hFFD7;
        rom[168][74] = 16'h001D;
        rom[168][75] = 16'h0016;
        rom[168][76] = 16'h0028;
        rom[168][77] = 16'hFFF4;
        rom[168][78] = 16'hFFCF;
        rom[168][79] = 16'h0007;
        rom[168][80] = 16'h001C;
        rom[168][81] = 16'h0025;
        rom[168][82] = 16'hFFE7;
        rom[168][83] = 16'hFFE1;
        rom[168][84] = 16'h0014;
        rom[168][85] = 16'h0006;
        rom[168][86] = 16'hFFBF;
        rom[168][87] = 16'h0038;
        rom[168][88] = 16'hFFF7;
        rom[168][89] = 16'hFFD0;
        rom[168][90] = 16'h0005;
        rom[168][91] = 16'h0002;
        rom[168][92] = 16'h001F;
        rom[168][93] = 16'hFFE4;
        rom[168][94] = 16'h0015;
        rom[168][95] = 16'hFFC2;
        rom[168][96] = 16'hFFBF;
        rom[168][97] = 16'h0032;
        rom[168][98] = 16'h0018;
        rom[168][99] = 16'h001B;
        rom[168][100] = 16'h0008;
        rom[168][101] = 16'hFFF9;
        rom[168][102] = 16'hFFFE;
        rom[168][103] = 16'h002B;
        rom[168][104] = 16'hFFC5;
        rom[168][105] = 16'h004D;
        rom[168][106] = 16'hFFEF;
        rom[168][107] = 16'h000D;
        rom[168][108] = 16'h0019;
        rom[168][109] = 16'hFFDF;
        rom[168][110] = 16'hFFEF;
        rom[168][111] = 16'h000F;
        rom[168][112] = 16'h0009;
        rom[168][113] = 16'h000C;
        rom[168][114] = 16'h002C;
        rom[168][115] = 16'h0020;
        rom[168][116] = 16'h0038;
        rom[168][117] = 16'hFFFE;
        rom[168][118] = 16'hFFFB;
        rom[168][119] = 16'hFFF5;
        rom[168][120] = 16'h001A;
        rom[168][121] = 16'h0011;
        rom[168][122] = 16'h0035;
        rom[168][123] = 16'hFFED;
        rom[168][124] = 16'h000C;
        rom[168][125] = 16'hFFFE;
        rom[168][126] = 16'h0006;
        rom[168][127] = 16'hFFD2;
        rom[169][0] = 16'h0011;
        rom[169][1] = 16'hFFE1;
        rom[169][2] = 16'hFFE1;
        rom[169][3] = 16'h0006;
        rom[169][4] = 16'hFFED;
        rom[169][5] = 16'hFFD8;
        rom[169][6] = 16'hFFF9;
        rom[169][7] = 16'hFFFD;
        rom[169][8] = 16'hFFEF;
        rom[169][9] = 16'h0018;
        rom[169][10] = 16'hFFF3;
        rom[169][11] = 16'h0025;
        rom[169][12] = 16'hFFB5;
        rom[169][13] = 16'h0012;
        rom[169][14] = 16'h0006;
        rom[169][15] = 16'hFFFE;
        rom[169][16] = 16'h0022;
        rom[169][17] = 16'h001A;
        rom[169][18] = 16'h001E;
        rom[169][19] = 16'hFFE9;
        rom[169][20] = 16'h003B;
        rom[169][21] = 16'h000C;
        rom[169][22] = 16'hFFCA;
        rom[169][23] = 16'h0038;
        rom[169][24] = 16'hFFF7;
        rom[169][25] = 16'h0016;
        rom[169][26] = 16'h001D;
        rom[169][27] = 16'h002D;
        rom[169][28] = 16'h0012;
        rom[169][29] = 16'h000A;
        rom[169][30] = 16'hFFDF;
        rom[169][31] = 16'h001C;
        rom[169][32] = 16'h0007;
        rom[169][33] = 16'h002C;
        rom[169][34] = 16'h0006;
        rom[169][35] = 16'h0009;
        rom[169][36] = 16'hFFF1;
        rom[169][37] = 16'h0001;
        rom[169][38] = 16'hFFF9;
        rom[169][39] = 16'h0044;
        rom[169][40] = 16'hFFB2;
        rom[169][41] = 16'h0030;
        rom[169][42] = 16'hFFEF;
        rom[169][43] = 16'hFFF4;
        rom[169][44] = 16'h0011;
        rom[169][45] = 16'h0005;
        rom[169][46] = 16'h0034;
        rom[169][47] = 16'h0057;
        rom[169][48] = 16'hFFC8;
        rom[169][49] = 16'hFFE1;
        rom[169][50] = 16'hFFC4;
        rom[169][51] = 16'hFFDD;
        rom[169][52] = 16'h0002;
        rom[169][53] = 16'h0020;
        rom[169][54] = 16'h001F;
        rom[169][55] = 16'hFFEA;
        rom[169][56] = 16'hFFD1;
        rom[169][57] = 16'h0026;
        rom[169][58] = 16'hFFED;
        rom[169][59] = 16'h0011;
        rom[169][60] = 16'hFFD8;
        rom[169][61] = 16'h0014;
        rom[169][62] = 16'hFFE1;
        rom[169][63] = 16'hFFFE;
        rom[169][64] = 16'hFFBA;
        rom[169][65] = 16'hFFF0;
        rom[169][66] = 16'hFFE1;
        rom[169][67] = 16'hFFE3;
        rom[169][68] = 16'hFFF7;
        rom[169][69] = 16'hFFF9;
        rom[169][70] = 16'h0005;
        rom[169][71] = 16'h0010;
        rom[169][72] = 16'h0011;
        rom[169][73] = 16'hFFBB;
        rom[169][74] = 16'h0019;
        rom[169][75] = 16'h0027;
        rom[169][76] = 16'hFFF5;
        rom[169][77] = 16'hFFDC;
        rom[169][78] = 16'hFFD9;
        rom[169][79] = 16'hFFEE;
        rom[169][80] = 16'hFFE4;
        rom[169][81] = 16'hFFFF;
        rom[169][82] = 16'hFFE2;
        rom[169][83] = 16'hFFED;
        rom[169][84] = 16'h0007;
        rom[169][85] = 16'hFFFE;
        rom[169][86] = 16'hFFFD;
        rom[169][87] = 16'hFFFA;
        rom[169][88] = 16'hFFF0;
        rom[169][89] = 16'h0024;
        rom[169][90] = 16'hFFD0;
        rom[169][91] = 16'h000B;
        rom[169][92] = 16'hFFF9;
        rom[169][93] = 16'h0002;
        rom[169][94] = 16'h0004;
        rom[169][95] = 16'hFFFE;
        rom[169][96] = 16'h0010;
        rom[169][97] = 16'h0012;
        rom[169][98] = 16'hFFDC;
        rom[169][99] = 16'hFFF7;
        rom[169][100] = 16'hFFF6;
        rom[169][101] = 16'hFFF5;
        rom[169][102] = 16'hFFD7;
        rom[169][103] = 16'h0026;
        rom[169][104] = 16'hFFD4;
        rom[169][105] = 16'h0022;
        rom[169][106] = 16'hFFDC;
        rom[169][107] = 16'h001E;
        rom[169][108] = 16'hFFFF;
        rom[169][109] = 16'hFFF3;
        rom[169][110] = 16'hFFDE;
        rom[169][111] = 16'h000C;
        rom[169][112] = 16'h0022;
        rom[169][113] = 16'hFFCD;
        rom[169][114] = 16'h0016;
        rom[169][115] = 16'hFFCF;
        rom[169][116] = 16'h0011;
        rom[169][117] = 16'h0011;
        rom[169][118] = 16'hFFD2;
        rom[169][119] = 16'hFFCD;
        rom[169][120] = 16'h000C;
        rom[169][121] = 16'h0015;
        rom[169][122] = 16'h0010;
        rom[169][123] = 16'hFFE7;
        rom[169][124] = 16'h0010;
        rom[169][125] = 16'hFFE4;
        rom[169][126] = 16'h0015;
        rom[169][127] = 16'h0011;
        rom[170][0] = 16'hFFE4;
        rom[170][1] = 16'h0010;
        rom[170][2] = 16'hFFE7;
        rom[170][3] = 16'h0029;
        rom[170][4] = 16'hFFF3;
        rom[170][5] = 16'h0011;
        rom[170][6] = 16'hFFFC;
        rom[170][7] = 16'h0012;
        rom[170][8] = 16'hFFF6;
        rom[170][9] = 16'h0002;
        rom[170][10] = 16'hFFD7;
        rom[170][11] = 16'hFFAA;
        rom[170][12] = 16'h0008;
        rom[170][13] = 16'hFFE7;
        rom[170][14] = 16'h0008;
        rom[170][15] = 16'hFFE2;
        rom[170][16] = 16'hFFFE;
        rom[170][17] = 16'h000C;
        rom[170][18] = 16'hFFDF;
        rom[170][19] = 16'hFFEE;
        rom[170][20] = 16'hFFAB;
        rom[170][21] = 16'hFFF2;
        rom[170][22] = 16'hFFFE;
        rom[170][23] = 16'h0026;
        rom[170][24] = 16'hFFF4;
        rom[170][25] = 16'h0018;
        rom[170][26] = 16'hFFEA;
        rom[170][27] = 16'h0002;
        rom[170][28] = 16'h002F;
        rom[170][29] = 16'hFFBC;
        rom[170][30] = 16'hFFE9;
        rom[170][31] = 16'hFFED;
        rom[170][32] = 16'hFFD4;
        rom[170][33] = 16'h0019;
        rom[170][34] = 16'h001B;
        rom[170][35] = 16'h001C;
        rom[170][36] = 16'hFFFA;
        rom[170][37] = 16'hFFEB;
        rom[170][38] = 16'hFFFE;
        rom[170][39] = 16'hFFB5;
        rom[170][40] = 16'h0010;
        rom[170][41] = 16'hFFD2;
        rom[170][42] = 16'h001D;
        rom[170][43] = 16'h001A;
        rom[170][44] = 16'hFFEF;
        rom[170][45] = 16'h0002;
        rom[170][46] = 16'h0016;
        rom[170][47] = 16'h001D;
        rom[170][48] = 16'hFFE9;
        rom[170][49] = 16'h0014;
        rom[170][50] = 16'h0008;
        rom[170][51] = 16'hFFE1;
        rom[170][52] = 16'h0003;
        rom[170][53] = 16'h0005;
        rom[170][54] = 16'hFFF9;
        rom[170][55] = 16'h002E;
        rom[170][56] = 16'hFFBC;
        rom[170][57] = 16'h0021;
        rom[170][58] = 16'hFFE1;
        rom[170][59] = 16'h000E;
        rom[170][60] = 16'h0002;
        rom[170][61] = 16'hFFDF;
        rom[170][62] = 16'h0011;
        rom[170][63] = 16'h0004;
        rom[170][64] = 16'hFFC6;
        rom[170][65] = 16'h0007;
        rom[170][66] = 16'h0010;
        rom[170][67] = 16'h0013;
        rom[170][68] = 16'h0008;
        rom[170][69] = 16'hFFFE;
        rom[170][70] = 16'h000C;
        rom[170][71] = 16'h0031;
        rom[170][72] = 16'hFFDD;
        rom[170][73] = 16'hFFEF;
        rom[170][74] = 16'h0001;
        rom[170][75] = 16'h0016;
        rom[170][76] = 16'hFFE1;
        rom[170][77] = 16'h000F;
        rom[170][78] = 16'hFFC3;
        rom[170][79] = 16'hFFF4;
        rom[170][80] = 16'h000D;
        rom[170][81] = 16'h0013;
        rom[170][82] = 16'h0018;
        rom[170][83] = 16'h0008;
        rom[170][84] = 16'hFFEB;
        rom[170][85] = 16'hFFFB;
        rom[170][86] = 16'hFFF4;
        rom[170][87] = 16'hFFEB;
        rom[170][88] = 16'hFFFB;
        rom[170][89] = 16'h0006;
        rom[170][90] = 16'h004D;
        rom[170][91] = 16'hFFCD;
        rom[170][92] = 16'hFFE4;
        rom[170][93] = 16'hFFE5;
        rom[170][94] = 16'hFFDE;
        rom[170][95] = 16'hFFFE;
        rom[170][96] = 16'hFFE5;
        rom[170][97] = 16'hFFDE;
        rom[170][98] = 16'hFFD2;
        rom[170][99] = 16'h001B;
        rom[170][100] = 16'h000F;
        rom[170][101] = 16'hFFE2;
        rom[170][102] = 16'h0029;
        rom[170][103] = 16'h000F;
        rom[170][104] = 16'hFFE2;
        rom[170][105] = 16'hFFD6;
        rom[170][106] = 16'h0007;
        rom[170][107] = 16'hFFF9;
        rom[170][108] = 16'hFFF7;
        rom[170][109] = 16'h000C;
        rom[170][110] = 16'hFFDE;
        rom[170][111] = 16'hFFFC;
        rom[170][112] = 16'hFFE3;
        rom[170][113] = 16'h0030;
        rom[170][114] = 16'hFFDF;
        rom[170][115] = 16'hFFFE;
        rom[170][116] = 16'h000A;
        rom[170][117] = 16'hFFE6;
        rom[170][118] = 16'hFFF0;
        rom[170][119] = 16'hFFF3;
        rom[170][120] = 16'hFFD0;
        rom[170][121] = 16'h0002;
        rom[170][122] = 16'hFFE5;
        rom[170][123] = 16'h0002;
        rom[170][124] = 16'hFFDC;
        rom[170][125] = 16'hFFFA;
        rom[170][126] = 16'h0029;
        rom[170][127] = 16'h0024;
        rom[171][0] = 16'h0008;
        rom[171][1] = 16'h0016;
        rom[171][2] = 16'hFFF0;
        rom[171][3] = 16'hFFC3;
        rom[171][4] = 16'h002E;
        rom[171][5] = 16'h000C;
        rom[171][6] = 16'h0026;
        rom[171][7] = 16'hFFFC;
        rom[171][8] = 16'hFFE5;
        rom[171][9] = 16'h0007;
        rom[171][10] = 16'h001D;
        rom[171][11] = 16'hFFF7;
        rom[171][12] = 16'hFFE0;
        rom[171][13] = 16'h001B;
        rom[171][14] = 16'hFFE9;
        rom[171][15] = 16'hFFDC;
        rom[171][16] = 16'h001B;
        rom[171][17] = 16'hFFF2;
        rom[171][18] = 16'h0013;
        rom[171][19] = 16'h002F;
        rom[171][20] = 16'h0002;
        rom[171][21] = 16'h0004;
        rom[171][22] = 16'h000A;
        rom[171][23] = 16'hFFEF;
        rom[171][24] = 16'h0011;
        rom[171][25] = 16'hFFF9;
        rom[171][26] = 16'hFFFD;
        rom[171][27] = 16'h0025;
        rom[171][28] = 16'hFFC6;
        rom[171][29] = 16'h0009;
        rom[171][30] = 16'h0040;
        rom[171][31] = 16'h000A;
        rom[171][32] = 16'h0008;
        rom[171][33] = 16'hFFE5;
        rom[171][34] = 16'hFFF9;
        rom[171][35] = 16'h000C;
        rom[171][36] = 16'h0012;
        rom[171][37] = 16'h004B;
        rom[171][38] = 16'h0026;
        rom[171][39] = 16'hFFFF;
        rom[171][40] = 16'hFFDC;
        rom[171][41] = 16'h002E;
        rom[171][42] = 16'hFFFE;
        rom[171][43] = 16'hFFC4;
        rom[171][44] = 16'h0004;
        rom[171][45] = 16'hFFFC;
        rom[171][46] = 16'h0015;
        rom[171][47] = 16'hFFD5;
        rom[171][48] = 16'hFFF3;
        rom[171][49] = 16'hFFE5;
        rom[171][50] = 16'hFFE1;
        rom[171][51] = 16'hFFDF;
        rom[171][52] = 16'hFFDC;
        rom[171][53] = 16'hFFD2;
        rom[171][54] = 16'h000D;
        rom[171][55] = 16'h002E;
        rom[171][56] = 16'h0008;
        rom[171][57] = 16'h0000;
        rom[171][58] = 16'hFFCF;
        rom[171][59] = 16'h0002;
        rom[171][60] = 16'h0002;
        rom[171][61] = 16'hFFFE;
        rom[171][62] = 16'hFFE4;
        rom[171][63] = 16'hFFFB;
        rom[171][64] = 16'hFFCB;
        rom[171][65] = 16'hFFF5;
        rom[171][66] = 16'hFFEA;
        rom[171][67] = 16'h0007;
        rom[171][68] = 16'hFFE6;
        rom[171][69] = 16'h001E;
        rom[171][70] = 16'h0002;
        rom[171][71] = 16'hFFC8;
        rom[171][72] = 16'h0018;
        rom[171][73] = 16'h000C;
        rom[171][74] = 16'hFFFF;
        rom[171][75] = 16'hFFF2;
        rom[171][76] = 16'hFFF8;
        rom[171][77] = 16'h0016;
        rom[171][78] = 16'hFFE7;
        rom[171][79] = 16'h0002;
        rom[171][80] = 16'h001E;
        rom[171][81] = 16'hFFFA;
        rom[171][82] = 16'h001B;
        rom[171][83] = 16'h001D;
        rom[171][84] = 16'h0002;
        rom[171][85] = 16'hFFF0;
        rom[171][86] = 16'h000C;
        rom[171][87] = 16'hFFE8;
        rom[171][88] = 16'hFFDE;
        rom[171][89] = 16'hFFD0;
        rom[171][90] = 16'hFFF4;
        rom[171][91] = 16'hFFEB;
        rom[171][92] = 16'hFFF8;
        rom[171][93] = 16'hFFBE;
        rom[171][94] = 16'hFFF6;
        rom[171][95] = 16'hFFD6;
        rom[171][96] = 16'hFFC8;
        rom[171][97] = 16'hFFD7;
        rom[171][98] = 16'h0006;
        rom[171][99] = 16'hFFE1;
        rom[171][100] = 16'hFFC9;
        rom[171][101] = 16'h002B;
        rom[171][102] = 16'hFFC3;
        rom[171][103] = 16'hFFEE;
        rom[171][104] = 16'hFFFE;
        rom[171][105] = 16'h0001;
        rom[171][106] = 16'hFFFE;
        rom[171][107] = 16'hFFF9;
        rom[171][108] = 16'hFFDF;
        rom[171][109] = 16'hFFDF;
        rom[171][110] = 16'hFFEA;
        rom[171][111] = 16'hFFF1;
        rom[171][112] = 16'h001B;
        rom[171][113] = 16'hFFEB;
        rom[171][114] = 16'hFFDF;
        rom[171][115] = 16'h0039;
        rom[171][116] = 16'h0007;
        rom[171][117] = 16'h0023;
        rom[171][118] = 16'hFFCD;
        rom[171][119] = 16'h0011;
        rom[171][120] = 16'h001B;
        rom[171][121] = 16'hFFD1;
        rom[171][122] = 16'h0013;
        rom[171][123] = 16'hFFF4;
        rom[171][124] = 16'hFFCB;
        rom[171][125] = 16'h0005;
        rom[171][126] = 16'hFFA6;
        rom[171][127] = 16'h0002;
        rom[172][0] = 16'h0011;
        rom[172][1] = 16'h0024;
        rom[172][2] = 16'hFFE5;
        rom[172][3] = 16'hFFFB;
        rom[172][4] = 16'h000A;
        rom[172][5] = 16'h0023;
        rom[172][6] = 16'h0010;
        rom[172][7] = 16'h0004;
        rom[172][8] = 16'h000D;
        rom[172][9] = 16'hFFDA;
        rom[172][10] = 16'h0011;
        rom[172][11] = 16'hFFD2;
        rom[172][12] = 16'h0007;
        rom[172][13] = 16'hFFFF;
        rom[172][14] = 16'hFFC2;
        rom[172][15] = 16'h0014;
        rom[172][16] = 16'h001F;
        rom[172][17] = 16'h0016;
        rom[172][18] = 16'hFFF8;
        rom[172][19] = 16'hFFFD;
        rom[172][20] = 16'hFFBC;
        rom[172][21] = 16'h0007;
        rom[172][22] = 16'hFFF5;
        rom[172][23] = 16'hFFEC;
        rom[172][24] = 16'hFFCD;
        rom[172][25] = 16'h0002;
        rom[172][26] = 16'h0021;
        rom[172][27] = 16'hFFF4;
        rom[172][28] = 16'hFFD1;
        rom[172][29] = 16'hFFE0;
        rom[172][30] = 16'h0016;
        rom[172][31] = 16'h001F;
        rom[172][32] = 16'hFFDE;
        rom[172][33] = 16'hFFF6;
        rom[172][34] = 16'h000F;
        rom[172][35] = 16'hFFDF;
        rom[172][36] = 16'h0039;
        rom[172][37] = 16'hFFF7;
        rom[172][38] = 16'hFFEF;
        rom[172][39] = 16'h000D;
        rom[172][40] = 16'h001F;
        rom[172][41] = 16'h0014;
        rom[172][42] = 16'hFFD4;
        rom[172][43] = 16'h0006;
        rom[172][44] = 16'h0003;
        rom[172][45] = 16'hFFC0;
        rom[172][46] = 16'hFFFF;
        rom[172][47] = 16'h001D;
        rom[172][48] = 16'h000D;
        rom[172][49] = 16'h0002;
        rom[172][50] = 16'hFFEF;
        rom[172][51] = 16'h0017;
        rom[172][52] = 16'hFFDC;
        rom[172][53] = 16'h0003;
        rom[172][54] = 16'h0014;
        rom[172][55] = 16'hFFE0;
        rom[172][56] = 16'h0022;
        rom[172][57] = 16'h000A;
        rom[172][58] = 16'h0011;
        rom[172][59] = 16'hFFE1;
        rom[172][60] = 16'h0025;
        rom[172][61] = 16'h000C;
        rom[172][62] = 16'h0000;
        rom[172][63] = 16'h001B;
        rom[172][64] = 16'h0011;
        rom[172][65] = 16'hFFE0;
        rom[172][66] = 16'h0016;
        rom[172][67] = 16'h002E;
        rom[172][68] = 16'h000B;
        rom[172][69] = 16'h0024;
        rom[172][70] = 16'h0000;
        rom[172][71] = 16'hFFB7;
        rom[172][72] = 16'hFFEA;
        rom[172][73] = 16'h0018;
        rom[172][74] = 16'h001C;
        rom[172][75] = 16'hFFD7;
        rom[172][76] = 16'hFFEE;
        rom[172][77] = 16'h0016;
        rom[172][78] = 16'hFFF7;
        rom[172][79] = 16'h0002;
        rom[172][80] = 16'hFFFF;
        rom[172][81] = 16'hFFF4;
        rom[172][82] = 16'h001C;
        rom[172][83] = 16'h0008;
        rom[172][84] = 16'hFFFA;
        rom[172][85] = 16'h0023;
        rom[172][86] = 16'h0024;
        rom[172][87] = 16'hFFD1;
        rom[172][88] = 16'h002C;
        rom[172][89] = 16'h0013;
        rom[172][90] = 16'hFFEE;
        rom[172][91] = 16'h0011;
        rom[172][92] = 16'hFFD7;
        rom[172][93] = 16'hFFFD;
        rom[172][94] = 16'hFFFF;
        rom[172][95] = 16'hFFEE;
        rom[172][96] = 16'h000F;
        rom[172][97] = 16'h0012;
        rom[172][98] = 16'h0024;
        rom[172][99] = 16'h000C;
        rom[172][100] = 16'hFFE7;
        rom[172][101] = 16'hFFED;
        rom[172][102] = 16'hFFEA;
        rom[172][103] = 16'h0002;
        rom[172][104] = 16'h0019;
        rom[172][105] = 16'h001B;
        rom[172][106] = 16'hFFF9;
        rom[172][107] = 16'hFFE4;
        rom[172][108] = 16'hFFDA;
        rom[172][109] = 16'hFFC4;
        rom[172][110] = 16'h0010;
        rom[172][111] = 16'h0021;
        rom[172][112] = 16'hFFC7;
        rom[172][113] = 16'h000C;
        rom[172][114] = 16'h0008;
        rom[172][115] = 16'hFFFE;
        rom[172][116] = 16'hFFE5;
        rom[172][117] = 16'h0001;
        rom[172][118] = 16'h0018;
        rom[172][119] = 16'h0016;
        rom[172][120] = 16'hFFFB;
        rom[172][121] = 16'h002A;
        rom[172][122] = 16'h000D;
        rom[172][123] = 16'hFFE1;
        rom[172][124] = 16'h000C;
        rom[172][125] = 16'h0005;
        rom[172][126] = 16'hFFCC;
        rom[172][127] = 16'hFFB8;
        rom[173][0] = 16'hFFFB;
        rom[173][1] = 16'hFFF6;
        rom[173][2] = 16'h0011;
        rom[173][3] = 16'hFFF1;
        rom[173][4] = 16'h0013;
        rom[173][5] = 16'h003F;
        rom[173][6] = 16'h0008;
        rom[173][7] = 16'hFFF4;
        rom[173][8] = 16'hFFF6;
        rom[173][9] = 16'h001E;
        rom[173][10] = 16'hFFF6;
        rom[173][11] = 16'h000C;
        rom[173][12] = 16'hFFEA;
        rom[173][13] = 16'h0024;
        rom[173][14] = 16'hFFD4;
        rom[173][15] = 16'h000B;
        rom[173][16] = 16'h0003;
        rom[173][17] = 16'hFFE1;
        rom[173][18] = 16'h0002;
        rom[173][19] = 16'hFFFD;
        rom[173][20] = 16'hFFEA;
        rom[173][21] = 16'hFFE5;
        rom[173][22] = 16'h0014;
        rom[173][23] = 16'hFFEB;
        rom[173][24] = 16'h0015;
        rom[173][25] = 16'h0008;
        rom[173][26] = 16'hFFEF;
        rom[173][27] = 16'h003C;
        rom[173][28] = 16'h0008;
        rom[173][29] = 16'h000E;
        rom[173][30] = 16'h0004;
        rom[173][31] = 16'h000D;
        rom[173][32] = 16'h0039;
        rom[173][33] = 16'hFFEA;
        rom[173][34] = 16'hFFF9;
        rom[173][35] = 16'h0034;
        rom[173][36] = 16'hFFDD;
        rom[173][37] = 16'hFFE2;
        rom[173][38] = 16'h001A;
        rom[173][39] = 16'hFFF9;
        rom[173][40] = 16'h001D;
        rom[173][41] = 16'h001A;
        rom[173][42] = 16'hFFA0;
        rom[173][43] = 16'hFFEB;
        rom[173][44] = 16'hFFFE;
        rom[173][45] = 16'h0017;
        rom[173][46] = 16'hFFFF;
        rom[173][47] = 16'hFFE9;
        rom[173][48] = 16'h0015;
        rom[173][49] = 16'h002C;
        rom[173][50] = 16'h0015;
        rom[173][51] = 16'hFFEF;
        rom[173][52] = 16'hFF97;
        rom[173][53] = 16'h0013;
        rom[173][54] = 16'h0017;
        rom[173][55] = 16'h0018;
        rom[173][56] = 16'hFFFE;
        rom[173][57] = 16'h0003;
        rom[173][58] = 16'hFFD3;
        rom[173][59] = 16'h0007;
        rom[173][60] = 16'hFFCB;
        rom[173][61] = 16'hFFF9;
        rom[173][62] = 16'h0033;
        rom[173][63] = 16'hFFE9;
        rom[173][64] = 16'hFFEA;
        rom[173][65] = 16'hFFF1;
        rom[173][66] = 16'h000C;
        rom[173][67] = 16'hFFDE;
        rom[173][68] = 16'hFFED;
        rom[173][69] = 16'hFFEB;
        rom[173][70] = 16'h0029;
        rom[173][71] = 16'hFFC2;
        rom[173][72] = 16'h000B;
        rom[173][73] = 16'h0006;
        rom[173][74] = 16'hFFCA;
        rom[173][75] = 16'hFFE3;
        rom[173][76] = 16'hFFEB;
        rom[173][77] = 16'hFFF6;
        rom[173][78] = 16'h000F;
        rom[173][79] = 16'h0012;
        rom[173][80] = 16'h0009;
        rom[173][81] = 16'hFFD1;
        rom[173][82] = 16'hFFF9;
        rom[173][83] = 16'h0007;
        rom[173][84] = 16'h0011;
        rom[173][85] = 16'h001B;
        rom[173][86] = 16'h001F;
        rom[173][87] = 16'hFFEA;
        rom[173][88] = 16'h001B;
        rom[173][89] = 16'h000B;
        rom[173][90] = 16'h0004;
        rom[173][91] = 16'hFFD8;
        rom[173][92] = 16'h0007;
        rom[173][93] = 16'hFFE5;
        rom[173][94] = 16'hFFE9;
        rom[173][95] = 16'h0029;
        rom[173][96] = 16'h0013;
        rom[173][97] = 16'h001C;
        rom[173][98] = 16'hFFEF;
        rom[173][99] = 16'hFFC6;
        rom[173][100] = 16'h0022;
        rom[173][101] = 16'h0007;
        rom[173][102] = 16'hFFE0;
        rom[173][103] = 16'hFFCF;
        rom[173][104] = 16'hFFEA;
        rom[173][105] = 16'hFFF1;
        rom[173][106] = 16'hFFEF;
        rom[173][107] = 16'hFFD4;
        rom[173][108] = 16'hFFFF;
        rom[173][109] = 16'hFFFB;
        rom[173][110] = 16'h0018;
        rom[173][111] = 16'h0000;
        rom[173][112] = 16'h0026;
        rom[173][113] = 16'h0027;
        rom[173][114] = 16'hFFD8;
        rom[173][115] = 16'hFFFE;
        rom[173][116] = 16'hFFED;
        rom[173][117] = 16'h001A;
        rom[173][118] = 16'h0005;
        rom[173][119] = 16'hFFFF;
        rom[173][120] = 16'hFFEE;
        rom[173][121] = 16'h0010;
        rom[173][122] = 16'h000C;
        rom[173][123] = 16'hFFCC;
        rom[173][124] = 16'h0017;
        rom[173][125] = 16'hFFF2;
        rom[173][126] = 16'hFFE7;
        rom[173][127] = 16'hFFB7;
        rom[174][0] = 16'hFFE0;
        rom[174][1] = 16'hFFEC;
        rom[174][2] = 16'h0016;
        rom[174][3] = 16'hFFF4;
        rom[174][4] = 16'h0028;
        rom[174][5] = 16'hFFF3;
        rom[174][6] = 16'hFFEC;
        rom[174][7] = 16'h000E;
        rom[174][8] = 16'hFFDE;
        rom[174][9] = 16'hFFC4;
        rom[174][10] = 16'hFFD7;
        rom[174][11] = 16'hFFE1;
        rom[174][12] = 16'h0025;
        rom[174][13] = 16'hFFD3;
        rom[174][14] = 16'hFFFA;
        rom[174][15] = 16'hFFF3;
        rom[174][16] = 16'h0012;
        rom[174][17] = 16'h0017;
        rom[174][18] = 16'hFFF9;
        rom[174][19] = 16'hFFF5;
        rom[174][20] = 16'h0017;
        rom[174][21] = 16'h0011;
        rom[174][22] = 16'h0013;
        rom[174][23] = 16'hFFCA;
        rom[174][24] = 16'hFFF6;
        rom[174][25] = 16'h0002;
        rom[174][26] = 16'h0009;
        rom[174][27] = 16'hFFEA;
        rom[174][28] = 16'h0001;
        rom[174][29] = 16'hFFE8;
        rom[174][30] = 16'h0019;
        rom[174][31] = 16'hFFFF;
        rom[174][32] = 16'hFFD5;
        rom[174][33] = 16'hFFF3;
        rom[174][34] = 16'hFFEF;
        rom[174][35] = 16'hFFEA;
        rom[174][36] = 16'h0006;
        rom[174][37] = 16'h001B;
        rom[174][38] = 16'hFFDC;
        rom[174][39] = 16'h0001;
        rom[174][40] = 16'hFFDA;
        rom[174][41] = 16'hFFE4;
        rom[174][42] = 16'hFFF8;
        rom[174][43] = 16'hFFFE;
        rom[174][44] = 16'h0005;
        rom[174][45] = 16'hFFEF;
        rom[174][46] = 16'h0003;
        rom[174][47] = 16'hFFEC;
        rom[174][48] = 16'h0010;
        rom[174][49] = 16'hFFDE;
        rom[174][50] = 16'h0007;
        rom[174][51] = 16'hFFD6;
        rom[174][52] = 16'h0012;
        rom[174][53] = 16'hFFF9;
        rom[174][54] = 16'h001E;
        rom[174][55] = 16'hFFED;
        rom[174][56] = 16'h0021;
        rom[174][57] = 16'hFFF8;
        rom[174][58] = 16'h0001;
        rom[174][59] = 16'h0011;
        rom[174][60] = 16'h0029;
        rom[174][61] = 16'h001F;
        rom[174][62] = 16'hFFF7;
        rom[174][63] = 16'hFFCA;
        rom[174][64] = 16'h000C;
        rom[174][65] = 16'h0003;
        rom[174][66] = 16'h0043;
        rom[174][67] = 16'hFFF5;
        rom[174][68] = 16'hFFEF;
        rom[174][69] = 16'hFFFE;
        rom[174][70] = 16'h001B;
        rom[174][71] = 16'h0016;
        rom[174][72] = 16'h003B;
        rom[174][73] = 16'hFFF4;
        rom[174][74] = 16'hFFE5;
        rom[174][75] = 16'h000A;
        rom[174][76] = 16'h0002;
        rom[174][77] = 16'h0008;
        rom[174][78] = 16'h001B;
        rom[174][79] = 16'hFFEF;
        rom[174][80] = 16'h0003;
        rom[174][81] = 16'h001F;
        rom[174][82] = 16'hFFF9;
        rom[174][83] = 16'hFFF6;
        rom[174][84] = 16'h000A;
        rom[174][85] = 16'hFFEF;
        rom[174][86] = 16'h000B;
        rom[174][87] = 16'h000C;
        rom[174][88] = 16'h001C;
        rom[174][89] = 16'hFFF5;
        rom[174][90] = 16'hFFFA;
        rom[174][91] = 16'h0002;
        rom[174][92] = 16'h0000;
        rom[174][93] = 16'hFFFF;
        rom[174][94] = 16'hFFEE;
        rom[174][95] = 16'hFFE6;
        rom[174][96] = 16'hFFDD;
        rom[174][97] = 16'hFFE3;
        rom[174][98] = 16'h0031;
        rom[174][99] = 16'h0045;
        rom[174][100] = 16'hFFEA;
        rom[174][101] = 16'h0024;
        rom[174][102] = 16'hFFF4;
        rom[174][103] = 16'h000C;
        rom[174][104] = 16'hFFE5;
        rom[174][105] = 16'hFFD4;
        rom[174][106] = 16'h0004;
        rom[174][107] = 16'hFFF3;
        rom[174][108] = 16'hFFF6;
        rom[174][109] = 16'hFFF0;
        rom[174][110] = 16'hFFF4;
        rom[174][111] = 16'h002A;
        rom[174][112] = 16'h0011;
        rom[174][113] = 16'h000A;
        rom[174][114] = 16'hFFFA;
        rom[174][115] = 16'h000B;
        rom[174][116] = 16'hFFF5;
        rom[174][117] = 16'hFFF4;
        rom[174][118] = 16'h0002;
        rom[174][119] = 16'h0032;
        rom[174][120] = 16'hFFFF;
        rom[174][121] = 16'hFFCC;
        rom[174][122] = 16'hFFFA;
        rom[174][123] = 16'hFFF5;
        rom[174][124] = 16'h0010;
        rom[174][125] = 16'h0001;
        rom[174][126] = 16'hFFFF;
        rom[174][127] = 16'h001B;
        rom[175][0] = 16'h0018;
        rom[175][1] = 16'h0023;
        rom[175][2] = 16'hFFFE;
        rom[175][3] = 16'hFF98;
        rom[175][4] = 16'h000F;
        rom[175][5] = 16'h001F;
        rom[175][6] = 16'hFFFD;
        rom[175][7] = 16'hFFFE;
        rom[175][8] = 16'hFFDF;
        rom[175][9] = 16'hFFEB;
        rom[175][10] = 16'hFFFF;
        rom[175][11] = 16'hFFF8;
        rom[175][12] = 16'hFFEF;
        rom[175][13] = 16'hFFFB;
        rom[175][14] = 16'hFFC4;
        rom[175][15] = 16'h001F;
        rom[175][16] = 16'h0003;
        rom[175][17] = 16'hFFEA;
        rom[175][18] = 16'h0034;
        rom[175][19] = 16'hFFFE;
        rom[175][20] = 16'h001C;
        rom[175][21] = 16'hFFF9;
        rom[175][22] = 16'hFFD1;
        rom[175][23] = 16'h0007;
        rom[175][24] = 16'h000B;
        rom[175][25] = 16'h001B;
        rom[175][26] = 16'hFFE9;
        rom[175][27] = 16'hFFE1;
        rom[175][28] = 16'h0006;
        rom[175][29] = 16'hFFE8;
        rom[175][30] = 16'h0011;
        rom[175][31] = 16'hFFC8;
        rom[175][32] = 16'h001B;
        rom[175][33] = 16'h001A;
        rom[175][34] = 16'hFFF2;
        rom[175][35] = 16'h001B;
        rom[175][36] = 16'h0005;
        rom[175][37] = 16'h0027;
        rom[175][38] = 16'hFFD4;
        rom[175][39] = 16'hFFEE;
        rom[175][40] = 16'hFFE7;
        rom[175][41] = 16'hFFC3;
        rom[175][42] = 16'hFFDF;
        rom[175][43] = 16'h0000;
        rom[175][44] = 16'h0007;
        rom[175][45] = 16'hFFF8;
        rom[175][46] = 16'hFFF4;
        rom[175][47] = 16'hFFFE;
        rom[175][48] = 16'h0007;
        rom[175][49] = 16'h0033;
        rom[175][50] = 16'hFFCF;
        rom[175][51] = 16'h0033;
        rom[175][52] = 16'hFFEA;
        rom[175][53] = 16'h0018;
        rom[175][54] = 16'hFFCE;
        rom[175][55] = 16'h0005;
        rom[175][56] = 16'h0035;
        rom[175][57] = 16'h000B;
        rom[175][58] = 16'hFFF2;
        rom[175][59] = 16'h0009;
        rom[175][60] = 16'h000D;
        rom[175][61] = 16'hFFC6;
        rom[175][62] = 16'hFFEA;
        rom[175][63] = 16'h0005;
        rom[175][64] = 16'hFFE8;
        rom[175][65] = 16'hFFFA;
        rom[175][66] = 16'h001B;
        rom[175][67] = 16'h001F;
        rom[175][68] = 16'h0020;
        rom[175][69] = 16'h0007;
        rom[175][70] = 16'hFFC9;
        rom[175][71] = 16'hFFDB;
        rom[175][72] = 16'hFFF1;
        rom[175][73] = 16'h0033;
        rom[175][74] = 16'hFFE9;
        rom[175][75] = 16'h0002;
        rom[175][76] = 16'hFFD8;
        rom[175][77] = 16'hFFCC;
        rom[175][78] = 16'hFFE9;
        rom[175][79] = 16'hFFC0;
        rom[175][80] = 16'hFFE0;
        rom[175][81] = 16'h000C;
        rom[175][82] = 16'hFFFE;
        rom[175][83] = 16'h0011;
        rom[175][84] = 16'h0008;
        rom[175][85] = 16'hFFDB;
        rom[175][86] = 16'h000D;
        rom[175][87] = 16'hFFE5;
        rom[175][88] = 16'h001F;
        rom[175][89] = 16'h0007;
        rom[175][90] = 16'hFFE6;
        rom[175][91] = 16'hFFF5;
        rom[175][92] = 16'h0011;
        rom[175][93] = 16'hFFFB;
        rom[175][94] = 16'hFFDB;
        rom[175][95] = 16'h0021;
        rom[175][96] = 16'hFFEE;
        rom[175][97] = 16'hFFEA;
        rom[175][98] = 16'h0008;
        rom[175][99] = 16'h0002;
        rom[175][100] = 16'h0003;
        rom[175][101] = 16'h001B;
        rom[175][102] = 16'h0005;
        rom[175][103] = 16'hFFFD;
        rom[175][104] = 16'h0003;
        rom[175][105] = 16'hFFE4;
        rom[175][106] = 16'hFFC5;
        rom[175][107] = 16'h001B;
        rom[175][108] = 16'h0000;
        rom[175][109] = 16'hFFFF;
        rom[175][110] = 16'h001D;
        rom[175][111] = 16'h0006;
        rom[175][112] = 16'h001B;
        rom[175][113] = 16'h0013;
        rom[175][114] = 16'h0038;
        rom[175][115] = 16'hFFF6;
        rom[175][116] = 16'hFFFD;
        rom[175][117] = 16'hFFD2;
        rom[175][118] = 16'h000B;
        rom[175][119] = 16'h0004;
        rom[175][120] = 16'h002E;
        rom[175][121] = 16'hFFFF;
        rom[175][122] = 16'h0005;
        rom[175][123] = 16'hFFF9;
        rom[175][124] = 16'hFFB3;
        rom[175][125] = 16'h000E;
        rom[175][126] = 16'hFFD2;
        rom[175][127] = 16'h0018;
        rom[176][0] = 16'h0012;
        rom[176][1] = 16'hFFF8;
        rom[176][2] = 16'h0025;
        rom[176][3] = 16'h001D;
        rom[176][4] = 16'hFFC5;
        rom[176][5] = 16'h0019;
        rom[176][6] = 16'h0006;
        rom[176][7] = 16'h000B;
        rom[176][8] = 16'hFFCC;
        rom[176][9] = 16'h0009;
        rom[176][10] = 16'hFFAD;
        rom[176][11] = 16'hFFE5;
        rom[176][12] = 16'hFFFE;
        rom[176][13] = 16'h0005;
        rom[176][14] = 16'hFFCF;
        rom[176][15] = 16'hFFE9;
        rom[176][16] = 16'hFFDD;
        rom[176][17] = 16'hFFF7;
        rom[176][18] = 16'hFFC6;
        rom[176][19] = 16'hFFF1;
        rom[176][20] = 16'hFFE5;
        rom[176][21] = 16'h0011;
        rom[176][22] = 16'hFFEE;
        rom[176][23] = 16'hFFAA;
        rom[176][24] = 16'h0029;
        rom[176][25] = 16'h002E;
        rom[176][26] = 16'hFFAF;
        rom[176][27] = 16'h0022;
        rom[176][28] = 16'hFFE8;
        rom[176][29] = 16'h0007;
        rom[176][30] = 16'hFFDC;
        rom[176][31] = 16'h001E;
        rom[176][32] = 16'hFFF9;
        rom[176][33] = 16'hFFDA;
        rom[176][34] = 16'h003F;
        rom[176][35] = 16'h0011;
        rom[176][36] = 16'hFFF4;
        rom[176][37] = 16'hFFC8;
        rom[176][38] = 16'h0016;
        rom[176][39] = 16'hFFC6;
        rom[176][40] = 16'hFFFE;
        rom[176][41] = 16'hFFE0;
        rom[176][42] = 16'hFFC2;
        rom[176][43] = 16'hFFCE;
        rom[176][44] = 16'h0012;
        rom[176][45] = 16'h0014;
        rom[176][46] = 16'hFFD4;
        rom[176][47] = 16'h0010;
        rom[176][48] = 16'hFFFF;
        rom[176][49] = 16'h0027;
        rom[176][50] = 16'h0012;
        rom[176][51] = 16'h000B;
        rom[176][52] = 16'h000C;
        rom[176][53] = 16'h0009;
        rom[176][54] = 16'h002E;
        rom[176][55] = 16'h002E;
        rom[176][56] = 16'hFFDE;
        rom[176][57] = 16'hFFE1;
        rom[176][58] = 16'hFFE5;
        rom[176][59] = 16'hFFDA;
        rom[176][60] = 16'h0006;
        rom[176][61] = 16'h000A;
        rom[176][62] = 16'h0002;
        rom[176][63] = 16'h000F;
        rom[176][64] = 16'h0000;
        rom[176][65] = 16'h0011;
        rom[176][66] = 16'hFFDF;
        rom[176][67] = 16'hFFB7;
        rom[176][68] = 16'h0002;
        rom[176][69] = 16'hFFFF;
        rom[176][70] = 16'h0028;
        rom[176][71] = 16'h0016;
        rom[176][72] = 16'h0011;
        rom[176][73] = 16'h0006;
        rom[176][74] = 16'h0004;
        rom[176][75] = 16'hFFDD;
        rom[176][76] = 16'h000B;
        rom[176][77] = 16'hFFCA;
        rom[176][78] = 16'hFFB8;
        rom[176][79] = 16'hFFDC;
        rom[176][80] = 16'h0013;
        rom[176][81] = 16'hFFF9;
        rom[176][82] = 16'hFFD3;
        rom[176][83] = 16'hFFEF;
        rom[176][84] = 16'h0009;
        rom[176][85] = 16'h0011;
        rom[176][86] = 16'hFFF4;
        rom[176][87] = 16'hFFFE;
        rom[176][88] = 16'h002E;
        rom[176][89] = 16'h0001;
        rom[176][90] = 16'hFFE0;
        rom[176][91] = 16'hFFFE;
        rom[176][92] = 16'hFFF9;
        rom[176][93] = 16'hFFD5;
        rom[176][94] = 16'h0016;
        rom[176][95] = 16'hFFB5;
        rom[176][96] = 16'hFFEA;
        rom[176][97] = 16'hFFFD;
        rom[176][98] = 16'h0017;
        rom[176][99] = 16'hFFF7;
        rom[176][100] = 16'h0006;
        rom[176][101] = 16'hFFF9;
        rom[176][102] = 16'h000F;
        rom[176][103] = 16'hFFEF;
        rom[176][104] = 16'h000C;
        rom[176][105] = 16'hFFDC;
        rom[176][106] = 16'h0000;
        rom[176][107] = 16'hFFE8;
        rom[176][108] = 16'h0020;
        rom[176][109] = 16'h0001;
        rom[176][110] = 16'h0002;
        rom[176][111] = 16'hFFB3;
        rom[176][112] = 16'hFFEE;
        rom[176][113] = 16'hFFC3;
        rom[176][114] = 16'h000A;
        rom[176][115] = 16'hFFFE;
        rom[176][116] = 16'hFFFD;
        rom[176][117] = 16'hFFD6;
        rom[176][118] = 16'h001F;
        rom[176][119] = 16'hFFF9;
        rom[176][120] = 16'h0008;
        rom[176][121] = 16'h0018;
        rom[176][122] = 16'hFFE5;
        rom[176][123] = 16'hFFFD;
        rom[176][124] = 16'h0007;
        rom[176][125] = 16'hFFD5;
        rom[176][126] = 16'h001E;
        rom[176][127] = 16'hFFDE;
        rom[177][0] = 16'h0020;
        rom[177][1] = 16'h0006;
        rom[177][2] = 16'h002D;
        rom[177][3] = 16'hFFE5;
        rom[177][4] = 16'hFFDB;
        rom[177][5] = 16'h0012;
        rom[177][6] = 16'h0002;
        rom[177][7] = 16'hFFD5;
        rom[177][8] = 16'hFFFE;
        rom[177][9] = 16'hFFEC;
        rom[177][10] = 16'hFFFB;
        rom[177][11] = 16'hFFBF;
        rom[177][12] = 16'h0001;
        rom[177][13] = 16'hFFFA;
        rom[177][14] = 16'hFFE6;
        rom[177][15] = 16'h0002;
        rom[177][16] = 16'hFFEF;
        rom[177][17] = 16'hFFD1;
        rom[177][18] = 16'hFFE1;
        rom[177][19] = 16'h0016;
        rom[177][20] = 16'hFFEA;
        rom[177][21] = 16'h001F;
        rom[177][22] = 16'h003A;
        rom[177][23] = 16'hFFC1;
        rom[177][24] = 16'hFFEA;
        rom[177][25] = 16'h002E;
        rom[177][26] = 16'hFFBF;
        rom[177][27] = 16'hFFEB;
        rom[177][28] = 16'hFFFD;
        rom[177][29] = 16'hFFE9;
        rom[177][30] = 16'hFFF9;
        rom[177][31] = 16'hFFF1;
        rom[177][32] = 16'h0007;
        rom[177][33] = 16'h000A;
        rom[177][34] = 16'h000C;
        rom[177][35] = 16'hFFD8;
        rom[177][36] = 16'hFFC6;
        rom[177][37] = 16'hFFE1;
        rom[177][38] = 16'hFFDD;
        rom[177][39] = 16'hFFE5;
        rom[177][40] = 16'h0005;
        rom[177][41] = 16'hFFCA;
        rom[177][42] = 16'h0038;
        rom[177][43] = 16'hFFC9;
        rom[177][44] = 16'hFFE5;
        rom[177][45] = 16'hFFE1;
        rom[177][46] = 16'hFFEE;
        rom[177][47] = 16'h0001;
        rom[177][48] = 16'hFFE8;
        rom[177][49] = 16'h002B;
        rom[177][50] = 16'h000F;
        rom[177][51] = 16'h002C;
        rom[177][52] = 16'h0002;
        rom[177][53] = 16'hFFD3;
        rom[177][54] = 16'hFFB0;
        rom[177][55] = 16'h001F;
        rom[177][56] = 16'h0002;
        rom[177][57] = 16'hFFF7;
        rom[177][58] = 16'hFFC0;
        rom[177][59] = 16'hFFB1;
        rom[177][60] = 16'h0018;
        rom[177][61] = 16'h0002;
        rom[177][62] = 16'hFFF2;
        rom[177][63] = 16'hFFA4;
        rom[177][64] = 16'hFFEC;
        rom[177][65] = 16'hFFD3;
        rom[177][66] = 16'hFFF9;
        rom[177][67] = 16'hFFFB;
        rom[177][68] = 16'h000A;
        rom[177][69] = 16'h0010;
        rom[177][70] = 16'h0013;
        rom[177][71] = 16'h0028;
        rom[177][72] = 16'hFFD9;
        rom[177][73] = 16'h0016;
        rom[177][74] = 16'hFFD9;
        rom[177][75] = 16'hFFF8;
        rom[177][76] = 16'hFFFB;
        rom[177][77] = 16'hFFD6;
        rom[177][78] = 16'hFFF9;
        rom[177][79] = 16'hFFAE;
        rom[177][80] = 16'h0023;
        rom[177][81] = 16'hFFEB;
        rom[177][82] = 16'hFFFD;
        rom[177][83] = 16'h000F;
        rom[177][84] = 16'h0024;
        rom[177][85] = 16'hFFF6;
        rom[177][86] = 16'hFFC7;
        rom[177][87] = 16'hFFEE;
        rom[177][88] = 16'h000A;
        rom[177][89] = 16'hFFE4;
        rom[177][90] = 16'h0028;
        rom[177][91] = 16'h0017;
        rom[177][92] = 16'h0011;
        rom[177][93] = 16'hFFFB;
        rom[177][94] = 16'hFFCE;
        rom[177][95] = 16'h0033;
        rom[177][96] = 16'hFFFE;
        rom[177][97] = 16'h0039;
        rom[177][98] = 16'h0018;
        rom[177][99] = 16'h0010;
        rom[177][100] = 16'hFFEE;
        rom[177][101] = 16'h0005;
        rom[177][102] = 16'h001F;
        rom[177][103] = 16'h0000;
        rom[177][104] = 16'h0021;
        rom[177][105] = 16'h0022;
        rom[177][106] = 16'hFFF6;
        rom[177][107] = 16'h0004;
        rom[177][108] = 16'h003E;
        rom[177][109] = 16'hFFE2;
        rom[177][110] = 16'hFFF9;
        rom[177][111] = 16'h0001;
        rom[177][112] = 16'h002F;
        rom[177][113] = 16'h0008;
        rom[177][114] = 16'h001B;
        rom[177][115] = 16'hFFEA;
        rom[177][116] = 16'h0003;
        rom[177][117] = 16'hFFE1;
        rom[177][118] = 16'hFFE5;
        rom[177][119] = 16'hFFE1;
        rom[177][120] = 16'h0023;
        rom[177][121] = 16'hFFD8;
        rom[177][122] = 16'h001D;
        rom[177][123] = 16'h0001;
        rom[177][124] = 16'hFFF8;
        rom[177][125] = 16'h0024;
        rom[177][126] = 16'h001C;
        rom[177][127] = 16'h0016;
        rom[178][0] = 16'h0005;
        rom[178][1] = 16'h0001;
        rom[178][2] = 16'h0008;
        rom[178][3] = 16'hFFFF;
        rom[178][4] = 16'h0015;
        rom[178][5] = 16'hFFD7;
        rom[178][6] = 16'hFFEF;
        rom[178][7] = 16'hFFED;
        rom[178][8] = 16'hFFD6;
        rom[178][9] = 16'h000B;
        rom[178][10] = 16'h0003;
        rom[178][11] = 16'h0007;
        rom[178][12] = 16'hFFE3;
        rom[178][13] = 16'hFFBF;
        rom[178][14] = 16'hFFE1;
        rom[178][15] = 16'h0004;
        rom[178][16] = 16'hFFF8;
        rom[178][17] = 16'hFFF3;
        rom[178][18] = 16'hFFDE;
        rom[178][19] = 16'h0001;
        rom[178][20] = 16'hFFF2;
        rom[178][21] = 16'hFFEC;
        rom[178][22] = 16'h0008;
        rom[178][23] = 16'h0011;
        rom[178][24] = 16'h0011;
        rom[178][25] = 16'hFFDC;
        rom[178][26] = 16'hFFED;
        rom[178][27] = 16'hFFF1;
        rom[178][28] = 16'h002C;
        rom[178][29] = 16'h000F;
        rom[178][30] = 16'hFFE2;
        rom[178][31] = 16'hFFE2;
        rom[178][32] = 16'hFFE6;
        rom[178][33] = 16'hFFE5;
        rom[178][34] = 16'h0023;
        rom[178][35] = 16'hFFDA;
        rom[178][36] = 16'hFFE1;
        rom[178][37] = 16'h002F;
        rom[178][38] = 16'h0002;
        rom[178][39] = 16'hFFED;
        rom[178][40] = 16'hFFDB;
        rom[178][41] = 16'hFFFA;
        rom[178][42] = 16'hFFE0;
        rom[178][43] = 16'hFFFC;
        rom[178][44] = 16'h000C;
        rom[178][45] = 16'hFFE6;
        rom[178][46] = 16'hFFF9;
        rom[178][47] = 16'hFFDC;
        rom[178][48] = 16'hFFE5;
        rom[178][49] = 16'hFFB5;
        rom[178][50] = 16'h0024;
        rom[178][51] = 16'h0011;
        rom[178][52] = 16'h0024;
        rom[178][53] = 16'hFFF4;
        rom[178][54] = 16'hFFAD;
        rom[178][55] = 16'hFFCD;
        rom[178][56] = 16'hFFFC;
        rom[178][57] = 16'h0009;
        rom[178][58] = 16'hFFF9;
        rom[178][59] = 16'h001B;
        rom[178][60] = 16'hFFF4;
        rom[178][61] = 16'hFFF5;
        rom[178][62] = 16'hFFB5;
        rom[178][63] = 16'hFFE1;
        rom[178][64] = 16'h001F;
        rom[178][65] = 16'hFFDB;
        rom[178][66] = 16'h0019;
        rom[178][67] = 16'h0018;
        rom[178][68] = 16'hFFBF;
        rom[178][69] = 16'hFFDE;
        rom[178][70] = 16'h001A;
        rom[178][71] = 16'h001B;
        rom[178][72] = 16'h000C;
        rom[178][73] = 16'hFFEC;
        rom[178][74] = 16'hFFCB;
        rom[178][75] = 16'h0018;
        rom[178][76] = 16'h0019;
        rom[178][77] = 16'hFFE5;
        rom[178][78] = 16'hFFEA;
        rom[178][79] = 16'hFFFE;
        rom[178][80] = 16'hFFBB;
        rom[178][81] = 16'hFFBA;
        rom[178][82] = 16'h0002;
        rom[178][83] = 16'hFFEE;
        rom[178][84] = 16'hFFF4;
        rom[178][85] = 16'hFFF5;
        rom[178][86] = 16'hFFE9;
        rom[178][87] = 16'h0036;
        rom[178][88] = 16'h0001;
        rom[178][89] = 16'hFFCE;
        rom[178][90] = 16'h0002;
        rom[178][91] = 16'hFFF1;
        rom[178][92] = 16'h0010;
        rom[178][93] = 16'hFFCE;
        rom[178][94] = 16'h0011;
        rom[178][95] = 16'hFFDD;
        rom[178][96] = 16'h0020;
        rom[178][97] = 16'hFFE7;
        rom[178][98] = 16'hFFE6;
        rom[178][99] = 16'hFFEC;
        rom[178][100] = 16'h001B;
        rom[178][101] = 16'h000C;
        rom[178][102] = 16'h0007;
        rom[178][103] = 16'h0016;
        rom[178][104] = 16'h0007;
        rom[178][105] = 16'hFFD9;
        rom[178][106] = 16'h0020;
        rom[178][107] = 16'h0006;
        rom[178][108] = 16'h000B;
        rom[178][109] = 16'h0019;
        rom[178][110] = 16'h0011;
        rom[178][111] = 16'hFFDC;
        rom[178][112] = 16'hFFD4;
        rom[178][113] = 16'hFFFE;
        rom[178][114] = 16'h0001;
        rom[178][115] = 16'hFFD9;
        rom[178][116] = 16'h0013;
        rom[178][117] = 16'h0010;
        rom[178][118] = 16'hFFE9;
        rom[178][119] = 16'h0015;
        rom[178][120] = 16'hFFF9;
        rom[178][121] = 16'h001B;
        rom[178][122] = 16'h0001;
        rom[178][123] = 16'h000C;
        rom[178][124] = 16'h0022;
        rom[178][125] = 16'h002E;
        rom[178][126] = 16'hFFEA;
        rom[178][127] = 16'h0001;
        rom[179][0] = 16'hFFF8;
        rom[179][1] = 16'hFFF9;
        rom[179][2] = 16'h0026;
        rom[179][3] = 16'hFFEC;
        rom[179][4] = 16'hFFC8;
        rom[179][5] = 16'hFFF2;
        rom[179][6] = 16'h0015;
        rom[179][7] = 16'h0002;
        rom[179][8] = 16'hFFF5;
        rom[179][9] = 16'h0023;
        rom[179][10] = 16'hFFF4;
        rom[179][11] = 16'hFFF2;
        rom[179][12] = 16'hFFEC;
        rom[179][13] = 16'hFFFE;
        rom[179][14] = 16'hFFEF;
        rom[179][15] = 16'h0016;
        rom[179][16] = 16'h0007;
        rom[179][17] = 16'h0002;
        rom[179][18] = 16'hFFEE;
        rom[179][19] = 16'hFFE7;
        rom[179][20] = 16'hFFFE;
        rom[179][21] = 16'h0011;
        rom[179][22] = 16'hFFAE;
        rom[179][23] = 16'hFFFE;
        rom[179][24] = 16'hFFED;
        rom[179][25] = 16'h0032;
        rom[179][26] = 16'h0006;
        rom[179][27] = 16'h0008;
        rom[179][28] = 16'hFFD9;
        rom[179][29] = 16'h0018;
        rom[179][30] = 16'hFFEA;
        rom[179][31] = 16'h0002;
        rom[179][32] = 16'hFFE5;
        rom[179][33] = 16'hFFFC;
        rom[179][34] = 16'h0005;
        rom[179][35] = 16'hFFFD;
        rom[179][36] = 16'h0002;
        rom[179][37] = 16'h001C;
        rom[179][38] = 16'hFFF3;
        rom[179][39] = 16'h0012;
        rom[179][40] = 16'h000B;
        rom[179][41] = 16'h0022;
        rom[179][42] = 16'hFFFB;
        rom[179][43] = 16'hFFFE;
        rom[179][44] = 16'h0021;
        rom[179][45] = 16'h0030;
        rom[179][46] = 16'hFFC3;
        rom[179][47] = 16'hFFE6;
        rom[179][48] = 16'h002F;
        rom[179][49] = 16'hFFE2;
        rom[179][50] = 16'h0009;
        rom[179][51] = 16'hFFD8;
        rom[179][52] = 16'h0006;
        rom[179][53] = 16'h001B;
        rom[179][54] = 16'hFFDC;
        rom[179][55] = 16'h0013;
        rom[179][56] = 16'h001C;
        rom[179][57] = 16'h0028;
        rom[179][58] = 16'h000B;
        rom[179][59] = 16'hFFCF;
        rom[179][60] = 16'hFFE1;
        rom[179][61] = 16'hFFD6;
        rom[179][62] = 16'hFFFA;
        rom[179][63] = 16'hFFF8;
        rom[179][64] = 16'h0001;
        rom[179][65] = 16'h0012;
        rom[179][66] = 16'hFFF7;
        rom[179][67] = 16'hFFCF;
        rom[179][68] = 16'h0014;
        rom[179][69] = 16'hFFDF;
        rom[179][70] = 16'hFFFD;
        rom[179][71] = 16'hFFFE;
        rom[179][72] = 16'h0016;
        rom[179][73] = 16'hFFD9;
        rom[179][74] = 16'h0016;
        rom[179][75] = 16'h0003;
        rom[179][76] = 16'h000C;
        rom[179][77] = 16'hFFE5;
        rom[179][78] = 16'hFFE9;
        rom[179][79] = 16'hFFFE;
        rom[179][80] = 16'h0015;
        rom[179][81] = 16'hFFE4;
        rom[179][82] = 16'hFFDF;
        rom[179][83] = 16'h0002;
        rom[179][84] = 16'hFFE8;
        rom[179][85] = 16'h0004;
        rom[179][86] = 16'h001D;
        rom[179][87] = 16'hFFF0;
        rom[179][88] = 16'hFFF9;
        rom[179][89] = 16'hFFDC;
        rom[179][90] = 16'hFFE0;
        rom[179][91] = 16'hFFF0;
        rom[179][92] = 16'hFFEA;
        rom[179][93] = 16'hFFAC;
        rom[179][94] = 16'h0018;
        rom[179][95] = 16'hFFDE;
        rom[179][96] = 16'h0011;
        rom[179][97] = 16'h001F;
        rom[179][98] = 16'hFFD9;
        rom[179][99] = 16'hFFCF;
        rom[179][100] = 16'h0001;
        rom[179][101] = 16'h0004;
        rom[179][102] = 16'hFFDB;
        rom[179][103] = 16'h0002;
        rom[179][104] = 16'hFFE5;
        rom[179][105] = 16'h0007;
        rom[179][106] = 16'h0018;
        rom[179][107] = 16'h0006;
        rom[179][108] = 16'hFFF0;
        rom[179][109] = 16'hFFE1;
        rom[179][110] = 16'hFFC3;
        rom[179][111] = 16'hFFF0;
        rom[179][112] = 16'hFFDC;
        rom[179][113] = 16'h0005;
        rom[179][114] = 16'hFFBB;
        rom[179][115] = 16'h0028;
        rom[179][116] = 16'hFFD8;
        rom[179][117] = 16'h001F;
        rom[179][118] = 16'hFFE5;
        rom[179][119] = 16'hFFE4;
        rom[179][120] = 16'h000E;
        rom[179][121] = 16'h0013;
        rom[179][122] = 16'hFFF1;
        rom[179][123] = 16'hFFB9;
        rom[179][124] = 16'hFFEF;
        rom[179][125] = 16'hFFE5;
        rom[179][126] = 16'hFFEF;
        rom[179][127] = 16'h000D;
        rom[180][0] = 16'hFFCF;
        rom[180][1] = 16'h0019;
        rom[180][2] = 16'hFFF9;
        rom[180][3] = 16'h0001;
        rom[180][4] = 16'hFFEA;
        rom[180][5] = 16'h0012;
        rom[180][6] = 16'hFFD8;
        rom[180][7] = 16'hFFF8;
        rom[180][8] = 16'h000D;
        rom[180][9] = 16'h0011;
        rom[180][10] = 16'h0007;
        rom[180][11] = 16'hFFEC;
        rom[180][12] = 16'h001A;
        rom[180][13] = 16'hFFF9;
        rom[180][14] = 16'h001C;
        rom[180][15] = 16'h0002;
        rom[180][16] = 16'hFFED;
        rom[180][17] = 16'hFFFC;
        rom[180][18] = 16'hFFF8;
        rom[180][19] = 16'hFFEF;
        rom[180][20] = 16'hFFC3;
        rom[180][21] = 16'hFFFE;
        rom[180][22] = 16'h0007;
        rom[180][23] = 16'h0010;
        rom[180][24] = 16'h001B;
        rom[180][25] = 16'hFFE7;
        rom[180][26] = 16'h0007;
        rom[180][27] = 16'hFFE5;
        rom[180][28] = 16'hFFE4;
        rom[180][29] = 16'h0017;
        rom[180][30] = 16'hFFF1;
        rom[180][31] = 16'hFFBD;
        rom[180][32] = 16'h0001;
        rom[180][33] = 16'h0004;
        rom[180][34] = 16'hFF9D;
        rom[180][35] = 16'hFFF6;
        rom[180][36] = 16'h0014;
        rom[180][37] = 16'hFFFE;
        rom[180][38] = 16'h0021;
        rom[180][39] = 16'hFFDB;
        rom[180][40] = 16'h001A;
        rom[180][41] = 16'hFFD7;
        rom[180][42] = 16'h0013;
        rom[180][43] = 16'hFFD6;
        rom[180][44] = 16'hFFF8;
        rom[180][45] = 16'h0018;
        rom[180][46] = 16'h0021;
        rom[180][47] = 16'h0039;
        rom[180][48] = 16'h001B;
        rom[180][49] = 16'h0007;
        rom[180][50] = 16'h001A;
        rom[180][51] = 16'hFFB9;
        rom[180][52] = 16'hFFAA;
        rom[180][53] = 16'hFFE6;
        rom[180][54] = 16'h000A;
        rom[180][55] = 16'hFFF0;
        rom[180][56] = 16'h0002;
        rom[180][57] = 16'hFFF3;
        rom[180][58] = 16'h0025;
        rom[180][59] = 16'h0032;
        rom[180][60] = 16'hFFE5;
        rom[180][61] = 16'hFFEC;
        rom[180][62] = 16'h000B;
        rom[180][63] = 16'hFFEA;
        rom[180][64] = 16'hFFDE;
        rom[180][65] = 16'h000F;
        rom[180][66] = 16'h0007;
        rom[180][67] = 16'hFFF9;
        rom[180][68] = 16'hFFEF;
        rom[180][69] = 16'h000A;
        rom[180][70] = 16'h0026;
        rom[180][71] = 16'hFFC0;
        rom[180][72] = 16'hFFE0;
        rom[180][73] = 16'h0004;
        rom[180][74] = 16'h0012;
        rom[180][75] = 16'h0002;
        rom[180][76] = 16'hFFE0;
        rom[180][77] = 16'h0026;
        rom[180][78] = 16'h0011;
        rom[180][79] = 16'h0012;
        rom[180][80] = 16'h0022;
        rom[180][81] = 16'h000C;
        rom[180][82] = 16'h0017;
        rom[180][83] = 16'h002C;
        rom[180][84] = 16'h0015;
        rom[180][85] = 16'hFFFF;
        rom[180][86] = 16'hFFF6;
        rom[180][87] = 16'hFFBF;
        rom[180][88] = 16'hFFD0;
        rom[180][89] = 16'h001A;
        rom[180][90] = 16'h0011;
        rom[180][91] = 16'hFFE8;
        rom[180][92] = 16'h0008;
        rom[180][93] = 16'h0033;
        rom[180][94] = 16'h0032;
        rom[180][95] = 16'hFFEF;
        rom[180][96] = 16'hFFFC;
        rom[180][97] = 16'hFFAF;
        rom[180][98] = 16'hFFF2;
        rom[180][99] = 16'h000A;
        rom[180][100] = 16'hFFB0;
        rom[180][101] = 16'hFFE2;
        rom[180][102] = 16'hFFF9;
        rom[180][103] = 16'h0002;
        rom[180][104] = 16'hFFE6;
        rom[180][105] = 16'hFFF1;
        rom[180][106] = 16'h000B;
        rom[180][107] = 16'hFFF9;
        rom[180][108] = 16'hFFBF;
        rom[180][109] = 16'h000E;
        rom[180][110] = 16'h000F;
        rom[180][111] = 16'hFFF1;
        rom[180][112] = 16'h0029;
        rom[180][113] = 16'h0000;
        rom[180][114] = 16'h0018;
        rom[180][115] = 16'hFFBE;
        rom[180][116] = 16'h0020;
        rom[180][117] = 16'h000F;
        rom[180][118] = 16'h0016;
        rom[180][119] = 16'h0011;
        rom[180][120] = 16'hFFEA;
        rom[180][121] = 16'hFFFE;
        rom[180][122] = 16'hFFFE;
        rom[180][123] = 16'h0016;
        rom[180][124] = 16'h000C;
        rom[180][125] = 16'hFFFE;
        rom[180][126] = 16'hFFC6;
        rom[180][127] = 16'hFFE6;
        rom[181][0] = 16'h0027;
        rom[181][1] = 16'hFFDB;
        rom[181][2] = 16'h0021;
        rom[181][3] = 16'hFFDB;
        rom[181][4] = 16'hFFDB;
        rom[181][5] = 16'h0017;
        rom[181][6] = 16'h0008;
        rom[181][7] = 16'h0005;
        rom[181][8] = 16'hFFF4;
        rom[181][9] = 16'h0008;
        rom[181][10] = 16'hFFFA;
        rom[181][11] = 16'hFFF2;
        rom[181][12] = 16'hFFFF;
        rom[181][13] = 16'hFFEA;
        rom[181][14] = 16'h000B;
        rom[181][15] = 16'h0006;
        rom[181][16] = 16'hFFD2;
        rom[181][17] = 16'hFFED;
        rom[181][18] = 16'h0022;
        rom[181][19] = 16'hFFEF;
        rom[181][20] = 16'hFFF7;
        rom[181][21] = 16'h0011;
        rom[181][22] = 16'h0006;
        rom[181][23] = 16'h0006;
        rom[181][24] = 16'h0017;
        rom[181][25] = 16'hFFFB;
        rom[181][26] = 16'hFFDF;
        rom[181][27] = 16'hFFE9;
        rom[181][28] = 16'hFFDF;
        rom[181][29] = 16'h000B;
        rom[181][30] = 16'hFFF5;
        rom[181][31] = 16'hFFFC;
        rom[181][32] = 16'h0015;
        rom[181][33] = 16'h0029;
        rom[181][34] = 16'hFFC8;
        rom[181][35] = 16'h000C;
        rom[181][36] = 16'hFFF7;
        rom[181][37] = 16'hFFE5;
        rom[181][38] = 16'h002E;
        rom[181][39] = 16'hFFEA;
        rom[181][40] = 16'hFFBA;
        rom[181][41] = 16'hFFDF;
        rom[181][42] = 16'hFFFA;
        rom[181][43] = 16'h0000;
        rom[181][44] = 16'hFFA0;
        rom[181][45] = 16'h0014;
        rom[181][46] = 16'h0011;
        rom[181][47] = 16'hFFDB;
        rom[181][48] = 16'h0002;
        rom[181][49] = 16'h001D;
        rom[181][50] = 16'h001F;
        rom[181][51] = 16'h001B;
        rom[181][52] = 16'h0007;
        rom[181][53] = 16'hFFEC;
        rom[181][54] = 16'h0029;
        rom[181][55] = 16'hFFDC;
        rom[181][56] = 16'h0016;
        rom[181][57] = 16'h0022;
        rom[181][58] = 16'h0016;
        rom[181][59] = 16'hFFEF;
        rom[181][60] = 16'hFFE6;
        rom[181][61] = 16'h0030;
        rom[181][62] = 16'hFFEB;
        rom[181][63] = 16'h0013;
        rom[181][64] = 16'h001E;
        rom[181][65] = 16'hFFEC;
        rom[181][66] = 16'hFFF1;
        rom[181][67] = 16'hFFEA;
        rom[181][68] = 16'hFFE7;
        rom[181][69] = 16'hFFF9;
        rom[181][70] = 16'h004D;
        rom[181][71] = 16'h000C;
        rom[181][72] = 16'h0029;
        rom[181][73] = 16'hFFE5;
        rom[181][74] = 16'hFFDE;
        rom[181][75] = 16'h0016;
        rom[181][76] = 16'h0004;
        rom[181][77] = 16'hFFD0;
        rom[181][78] = 16'hFFFE;
        rom[181][79] = 16'hFFD7;
        rom[181][80] = 16'hFFFE;
        rom[181][81] = 16'h0033;
        rom[181][82] = 16'hFFEB;
        rom[181][83] = 16'hFFF5;
        rom[181][84] = 16'h0007;
        rom[181][85] = 16'hFFF2;
        rom[181][86] = 16'h0001;
        rom[181][87] = 16'hFFF1;
        rom[181][88] = 16'h0011;
        rom[181][89] = 16'h0033;
        rom[181][90] = 16'hFFF5;
        rom[181][91] = 16'hFFB8;
        rom[181][92] = 16'hFFCD;
        rom[181][93] = 16'h000F;
        rom[181][94] = 16'hFFB3;
        rom[181][95] = 16'h0002;
        rom[181][96] = 16'hFFF0;
        rom[181][97] = 16'h0001;
        rom[181][98] = 16'hFFF5;
        rom[181][99] = 16'h0011;
        rom[181][100] = 16'hFFE8;
        rom[181][101] = 16'h001C;
        rom[181][102] = 16'hFFEA;
        rom[181][103] = 16'h000E;
        rom[181][104] = 16'hFFF5;
        rom[181][105] = 16'hFFAB;
        rom[181][106] = 16'hFFFB;
        rom[181][107] = 16'h0012;
        rom[181][108] = 16'h001F;
        rom[181][109] = 16'h001D;
        rom[181][110] = 16'hFFF2;
        rom[181][111] = 16'hFFEE;
        rom[181][112] = 16'hFFF8;
        rom[181][113] = 16'hFFFC;
        rom[181][114] = 16'hFFFE;
        rom[181][115] = 16'hFFC1;
        rom[181][116] = 16'h0002;
        rom[181][117] = 16'hFFE7;
        rom[181][118] = 16'h0001;
        rom[181][119] = 16'h001E;
        rom[181][120] = 16'h0013;
        rom[181][121] = 16'hFFFA;
        rom[181][122] = 16'h0006;
        rom[181][123] = 16'hFFF7;
        rom[181][124] = 16'hFFE5;
        rom[181][125] = 16'h0001;
        rom[181][126] = 16'hFFE8;
        rom[181][127] = 16'hFFF0;
        rom[182][0] = 16'h0005;
        rom[182][1] = 16'hFFC3;
        rom[182][2] = 16'hFFFB;
        rom[182][3] = 16'h0030;
        rom[182][4] = 16'hFFF9;
        rom[182][5] = 16'hFFC7;
        rom[182][6] = 16'hFFD7;
        rom[182][7] = 16'hFFF6;
        rom[182][8] = 16'hFFD2;
        rom[182][9] = 16'h001F;
        rom[182][10] = 16'hFFFD;
        rom[182][11] = 16'h002E;
        rom[182][12] = 16'hFFE0;
        rom[182][13] = 16'h0007;
        rom[182][14] = 16'hFFE6;
        rom[182][15] = 16'h0011;
        rom[182][16] = 16'hFFF4;
        rom[182][17] = 16'hFFF0;
        rom[182][18] = 16'h004F;
        rom[182][19] = 16'hFFF4;
        rom[182][20] = 16'h0044;
        rom[182][21] = 16'h000A;
        rom[182][22] = 16'h0024;
        rom[182][23] = 16'h0006;
        rom[182][24] = 16'hFFFC;
        rom[182][25] = 16'h0010;
        rom[182][26] = 16'h0008;
        rom[182][27] = 16'hFFF6;
        rom[182][28] = 16'hFFF4;
        rom[182][29] = 16'hFFEC;
        rom[182][30] = 16'h0003;
        rom[182][31] = 16'hFFF1;
        rom[182][32] = 16'hFFF5;
        rom[182][33] = 16'h001B;
        rom[182][34] = 16'hFFF3;
        rom[182][35] = 16'hFFFA;
        rom[182][36] = 16'hFFDC;
        rom[182][37] = 16'hFFE5;
        rom[182][38] = 16'h0021;
        rom[182][39] = 16'hFFBB;
        rom[182][40] = 16'hFFEF;
        rom[182][41] = 16'hFFDE;
        rom[182][42] = 16'h0024;
        rom[182][43] = 16'hFFCC;
        rom[182][44] = 16'hFFDC;
        rom[182][45] = 16'h0000;
        rom[182][46] = 16'h0012;
        rom[182][47] = 16'hFFE3;
        rom[182][48] = 16'hFFE1;
        rom[182][49] = 16'hFFDE;
        rom[182][50] = 16'hFFCE;
        rom[182][51] = 16'h0002;
        rom[182][52] = 16'h0008;
        rom[182][53] = 16'hFFF4;
        rom[182][54] = 16'hFFE6;
        rom[182][55] = 16'h0023;
        rom[182][56] = 16'h0007;
        rom[182][57] = 16'hFFF3;
        rom[182][58] = 16'h0017;
        rom[182][59] = 16'hFFFA;
        rom[182][60] = 16'hFFAD;
        rom[182][61] = 16'hFFCA;
        rom[182][62] = 16'hFFF6;
        rom[182][63] = 16'hFFB9;
        rom[182][64] = 16'h000D;
        rom[182][65] = 16'h000C;
        rom[182][66] = 16'hFFD2;
        rom[182][67] = 16'hFFF7;
        rom[182][68] = 16'hFFE9;
        rom[182][69] = 16'hFFEA;
        rom[182][70] = 16'hFFF6;
        rom[182][71] = 16'hFFF4;
        rom[182][72] = 16'hFFF2;
        rom[182][73] = 16'hFFFC;
        rom[182][74] = 16'hFFD7;
        rom[182][75] = 16'h0000;
        rom[182][76] = 16'h001E;
        rom[182][77] = 16'hFFF4;
        rom[182][78] = 16'hFFD5;
        rom[182][79] = 16'hFFED;
        rom[182][80] = 16'hFFAC;
        rom[182][81] = 16'hFFE6;
        rom[182][82] = 16'hFFEF;
        rom[182][83] = 16'h0002;
        rom[182][84] = 16'hFFE1;
        rom[182][85] = 16'h000E;
        rom[182][86] = 16'h000A;
        rom[182][87] = 16'h0019;
        rom[182][88] = 16'h0030;
        rom[182][89] = 16'hFFFB;
        rom[182][90] = 16'h002A;
        rom[182][91] = 16'h0011;
        rom[182][92] = 16'h0021;
        rom[182][93] = 16'hFFE8;
        rom[182][94] = 16'hFFE3;
        rom[182][95] = 16'h001B;
        rom[182][96] = 16'hFFEF;
        rom[182][97] = 16'hFFEA;
        rom[182][98] = 16'hFFD0;
        rom[182][99] = 16'hFFD8;
        rom[182][100] = 16'hFFDC;
        rom[182][101] = 16'hFFFF;
        rom[182][102] = 16'h0010;
        rom[182][103] = 16'hFFEF;
        rom[182][104] = 16'h0027;
        rom[182][105] = 16'hFFFA;
        rom[182][106] = 16'hFFEF;
        rom[182][107] = 16'h001A;
        rom[182][108] = 16'hFFEA;
        rom[182][109] = 16'hFFF4;
        rom[182][110] = 16'hFFE7;
        rom[182][111] = 16'hFFDD;
        rom[182][112] = 16'h0002;
        rom[182][113] = 16'h0025;
        rom[182][114] = 16'hFFDE;
        rom[182][115] = 16'h001F;
        rom[182][116] = 16'h0011;
        rom[182][117] = 16'hFFFA;
        rom[182][118] = 16'hFFBA;
        rom[182][119] = 16'hFFE4;
        rom[182][120] = 16'h0002;
        rom[182][121] = 16'h0003;
        rom[182][122] = 16'h001C;
        rom[182][123] = 16'h001D;
        rom[182][124] = 16'hFFFE;
        rom[182][125] = 16'h0002;
        rom[182][126] = 16'h0010;
        rom[182][127] = 16'h001D;
        rom[183][0] = 16'h0002;
        rom[183][1] = 16'h000F;
        rom[183][2] = 16'h0006;
        rom[183][3] = 16'hFFD1;
        rom[183][4] = 16'hFFD6;
        rom[183][5] = 16'h0019;
        rom[183][6] = 16'hFFBF;
        rom[183][7] = 16'h0007;
        rom[183][8] = 16'h0009;
        rom[183][9] = 16'h0033;
        rom[183][10] = 16'h0009;
        rom[183][11] = 16'hFFF3;
        rom[183][12] = 16'h0031;
        rom[183][13] = 16'hFFEF;
        rom[183][14] = 16'hFFED;
        rom[183][15] = 16'h0009;
        rom[183][16] = 16'h0007;
        rom[183][17] = 16'hFFE9;
        rom[183][18] = 16'h000D;
        rom[183][19] = 16'h0010;
        rom[183][20] = 16'hFFEA;
        rom[183][21] = 16'hFFF9;
        rom[183][22] = 16'hFFEE;
        rom[183][23] = 16'h0009;
        rom[183][24] = 16'h001D;
        rom[183][25] = 16'h0014;
        rom[183][26] = 16'h0011;
        rom[183][27] = 16'hFFDC;
        rom[183][28] = 16'hFFB5;
        rom[183][29] = 16'hFFCB;
        rom[183][30] = 16'hFFEA;
        rom[183][31] = 16'hFFF1;
        rom[183][32] = 16'hFFE8;
        rom[183][33] = 16'h000B;
        rom[183][34] = 16'hFFC6;
        rom[183][35] = 16'hFFF8;
        rom[183][36] = 16'h0009;
        rom[183][37] = 16'hFFFB;
        rom[183][38] = 16'h0033;
        rom[183][39] = 16'hFFEF;
        rom[183][40] = 16'hFFDB;
        rom[183][41] = 16'hFFF9;
        rom[183][42] = 16'h001A;
        rom[183][43] = 16'h0006;
        rom[183][44] = 16'hFFE6;
        rom[183][45] = 16'h0012;
        rom[183][46] = 16'h0007;
        rom[183][47] = 16'h0026;
        rom[183][48] = 16'h001F;
        rom[183][49] = 16'h002C;
        rom[183][50] = 16'h0009;
        rom[183][51] = 16'hFFC7;
        rom[183][52] = 16'hFFD6;
        rom[183][53] = 16'hFFE5;
        rom[183][54] = 16'hFFD4;
        rom[183][55] = 16'h0011;
        rom[183][56] = 16'hFFFD;
        rom[183][57] = 16'h000E;
        rom[183][58] = 16'h0011;
        rom[183][59] = 16'hFFE7;
        rom[183][60] = 16'h0001;
        rom[183][61] = 16'hFFE2;
        rom[183][62] = 16'h0003;
        rom[183][63] = 16'h0012;
        rom[183][64] = 16'hFFC2;
        rom[183][65] = 16'hFFF8;
        rom[183][66] = 16'hFFFF;
        rom[183][67] = 16'h001B;
        rom[183][68] = 16'hFFD7;
        rom[183][69] = 16'h0012;
        rom[183][70] = 16'h0020;
        rom[183][71] = 16'hFFBF;
        rom[183][72] = 16'h000A;
        rom[183][73] = 16'hFFF3;
        rom[183][74] = 16'h0008;
        rom[183][75] = 16'h0010;
        rom[183][76] = 16'h000F;
        rom[183][77] = 16'hFFF2;
        rom[183][78] = 16'hFFE1;
        rom[183][79] = 16'hFFFE;
        rom[183][80] = 16'h002F;
        rom[183][81] = 16'hFFF4;
        rom[183][82] = 16'h001C;
        rom[183][83] = 16'h0018;
        rom[183][84] = 16'hFFF9;
        rom[183][85] = 16'h001A;
        rom[183][86] = 16'hFFFB;
        rom[183][87] = 16'hFFCB;
        rom[183][88] = 16'hFFDB;
        rom[183][89] = 16'hFFE2;
        rom[183][90] = 16'hFFFC;
        rom[183][91] = 16'h0007;
        rom[183][92] = 16'hFFE5;
        rom[183][93] = 16'hFFDA;
        rom[183][94] = 16'hFFDC;
        rom[183][95] = 16'hFFC4;
        rom[183][96] = 16'hFFD7;
        rom[183][97] = 16'h0006;
        rom[183][98] = 16'hFFE0;
        rom[183][99] = 16'h0024;
        rom[183][100] = 16'hFFC4;
        rom[183][101] = 16'hFFDD;
        rom[183][102] = 16'hFFDB;
        rom[183][103] = 16'hFFCD;
        rom[183][104] = 16'hFFE0;
        rom[183][105] = 16'hFFD7;
        rom[183][106] = 16'hFFF5;
        rom[183][107] = 16'h0022;
        rom[183][108] = 16'hFFC4;
        rom[183][109] = 16'hFFF6;
        rom[183][110] = 16'h0018;
        rom[183][111] = 16'h0007;
        rom[183][112] = 16'hFFA3;
        rom[183][113] = 16'h002E;
        rom[183][114] = 16'hFFE7;
        rom[183][115] = 16'hFFDF;
        rom[183][116] = 16'hFFFE;
        rom[183][117] = 16'h0022;
        rom[183][118] = 16'h0020;
        rom[183][119] = 16'h002D;
        rom[183][120] = 16'hFFE1;
        rom[183][121] = 16'h000E;
        rom[183][122] = 16'hFFDE;
        rom[183][123] = 16'h0011;
        rom[183][124] = 16'hFFCD;
        rom[183][125] = 16'hFFEA;
        rom[183][126] = 16'hFFEB;
        rom[183][127] = 16'h0022;
        rom[184][0] = 16'h000C;
        rom[184][1] = 16'h0016;
        rom[184][2] = 16'hFFE6;
        rom[184][3] = 16'hFFF4;
        rom[184][4] = 16'hFFEF;
        rom[184][5] = 16'hFFFD;
        rom[184][6] = 16'hFFF6;
        rom[184][7] = 16'h0010;
        rom[184][8] = 16'h001A;
        rom[184][9] = 16'hFFE2;
        rom[184][10] = 16'hFFCB;
        rom[184][11] = 16'hFFC7;
        rom[184][12] = 16'h0011;
        rom[184][13] = 16'h0012;
        rom[184][14] = 16'h0016;
        rom[184][15] = 16'hFFF5;
        rom[184][16] = 16'h000F;
        rom[184][17] = 16'hFFC0;
        rom[184][18] = 16'hFFF9;
        rom[184][19] = 16'hFFEF;
        rom[184][20] = 16'hFFDE;
        rom[184][21] = 16'h0028;
        rom[184][22] = 16'hFFCF;
        rom[184][23] = 16'hFFD2;
        rom[184][24] = 16'h000C;
        rom[184][25] = 16'h0034;
        rom[184][26] = 16'h0002;
        rom[184][27] = 16'hFFC8;
        rom[184][28] = 16'hFFB1;
        rom[184][29] = 16'hFFD7;
        rom[184][30] = 16'h0007;
        rom[184][31] = 16'h0029;
        rom[184][32] = 16'hFFA7;
        rom[184][33] = 16'h0026;
        rom[184][34] = 16'hFFEE;
        rom[184][35] = 16'hFFD7;
        rom[184][36] = 16'h0011;
        rom[184][37] = 16'hFFE5;
        rom[184][38] = 16'h0007;
        rom[184][39] = 16'hFFD8;
        rom[184][40] = 16'hFFE7;
        rom[184][41] = 16'h000E;
        rom[184][42] = 16'h002F;
        rom[184][43] = 16'h0024;
        rom[184][44] = 16'hFFE3;
        rom[184][45] = 16'hFFE3;
        rom[184][46] = 16'h0026;
        rom[184][47] = 16'h0016;
        rom[184][48] = 16'h0011;
        rom[184][49] = 16'h0002;
        rom[184][50] = 16'hFFFB;
        rom[184][51] = 16'hFFCE;
        rom[184][52] = 16'hFFF9;
        rom[184][53] = 16'hFFC9;
        rom[184][54] = 16'h0018;
        rom[184][55] = 16'hFFF3;
        rom[184][56] = 16'hFFE6;
        rom[184][57] = 16'h0005;
        rom[184][58] = 16'h0049;
        rom[184][59] = 16'hFFD0;
        rom[184][60] = 16'h0011;
        rom[184][61] = 16'hFFF4;
        rom[184][62] = 16'h0014;
        rom[184][63] = 16'h0002;
        rom[184][64] = 16'h0012;
        rom[184][65] = 16'h0002;
        rom[184][66] = 16'hFFD5;
        rom[184][67] = 16'hFFE7;
        rom[184][68] = 16'hFFFC;
        rom[184][69] = 16'hFFEA;
        rom[184][70] = 16'hFFFF;
        rom[184][71] = 16'h0019;
        rom[184][72] = 16'h000F;
        rom[184][73] = 16'hFFD7;
        rom[184][74] = 16'h0015;
        rom[184][75] = 16'h0018;
        rom[184][76] = 16'h0011;
        rom[184][77] = 16'hFFE4;
        rom[184][78] = 16'hFFE0;
        rom[184][79] = 16'h004F;
        rom[184][80] = 16'hFFF5;
        rom[184][81] = 16'h0018;
        rom[184][82] = 16'h0004;
        rom[184][83] = 16'hFFFE;
        rom[184][84] = 16'h000E;
        rom[184][85] = 16'hFFDC;
        rom[184][86] = 16'h0015;
        rom[184][87] = 16'hFFF6;
        rom[184][88] = 16'h002C;
        rom[184][89] = 16'hFFC3;
        rom[184][90] = 16'h0013;
        rom[184][91] = 16'h001B;
        rom[184][92] = 16'hFFFD;
        rom[184][93] = 16'hFFCD;
        rom[184][94] = 16'hFFE6;
        rom[184][95] = 16'hFFBF;
        rom[184][96] = 16'hFFDF;
        rom[184][97] = 16'hFFDD;
        rom[184][98] = 16'h0029;
        rom[184][99] = 16'h0018;
        rom[184][100] = 16'hFFDC;
        rom[184][101] = 16'h000A;
        rom[184][102] = 16'h0029;
        rom[184][103] = 16'hFFE1;
        rom[184][104] = 16'h001B;
        rom[184][105] = 16'h000C;
        rom[184][106] = 16'hFFF3;
        rom[184][107] = 16'h0009;
        rom[184][108] = 16'hFFE1;
        rom[184][109] = 16'hFFD9;
        rom[184][110] = 16'h0002;
        rom[184][111] = 16'hFFFE;
        rom[184][112] = 16'hFFE5;
        rom[184][113] = 16'h0027;
        rom[184][114] = 16'hFFDC;
        rom[184][115] = 16'h0014;
        rom[184][116] = 16'hFFEF;
        rom[184][117] = 16'hFFF4;
        rom[184][118] = 16'hFFFF;
        rom[184][119] = 16'h0009;
        rom[184][120] = 16'h0015;
        rom[184][121] = 16'hFFCF;
        rom[184][122] = 16'hFFE5;
        rom[184][123] = 16'h0007;
        rom[184][124] = 16'hFFF1;
        rom[184][125] = 16'hFFFF;
        rom[184][126] = 16'hFFD2;
        rom[184][127] = 16'h0006;
        rom[185][0] = 16'h0037;
        rom[185][1] = 16'hFFE0;
        rom[185][2] = 16'hFFF9;
        rom[185][3] = 16'hFFF2;
        rom[185][4] = 16'hFFF4;
        rom[185][5] = 16'hFFD9;
        rom[185][6] = 16'h0002;
        rom[185][7] = 16'hFFFD;
        rom[185][8] = 16'hFFF7;
        rom[185][9] = 16'h001B;
        rom[185][10] = 16'h0017;
        rom[185][11] = 16'h001D;
        rom[185][12] = 16'hFFCA;
        rom[185][13] = 16'hFFE3;
        rom[185][14] = 16'hFFE5;
        rom[185][15] = 16'hFFED;
        rom[185][16] = 16'hFFEF;
        rom[185][17] = 16'hFFFE;
        rom[185][18] = 16'hFFF8;
        rom[185][19] = 16'h0017;
        rom[185][20] = 16'h000C;
        rom[185][21] = 16'h0015;
        rom[185][22] = 16'h0008;
        rom[185][23] = 16'h000C;
        rom[185][24] = 16'h0009;
        rom[185][25] = 16'hFFD8;
        rom[185][26] = 16'hFFE7;
        rom[185][27] = 16'hFFEA;
        rom[185][28] = 16'hFFDA;
        rom[185][29] = 16'hFFD7;
        rom[185][30] = 16'hFFEC;
        rom[185][31] = 16'hFFF7;
        rom[185][32] = 16'hFFF0;
        rom[185][33] = 16'h0007;
        rom[185][34] = 16'hFFF0;
        rom[185][35] = 16'hFFF4;
        rom[185][36] = 16'hFFE3;
        rom[185][37] = 16'hFFDC;
        rom[185][38] = 16'h001F;
        rom[185][39] = 16'h0029;
        rom[185][40] = 16'hFFD0;
        rom[185][41] = 16'h0014;
        rom[185][42] = 16'hFFC7;
        rom[185][43] = 16'h0017;
        rom[185][44] = 16'h000C;
        rom[185][45] = 16'h0011;
        rom[185][46] = 16'hFFD9;
        rom[185][47] = 16'hFFE6;
        rom[185][48] = 16'hFFDB;
        rom[185][49] = 16'hFFE6;
        rom[185][50] = 16'h000C;
        rom[185][51] = 16'h0029;
        rom[185][52] = 16'h0007;
        rom[185][53] = 16'hFFEF;
        rom[185][54] = 16'h000B;
        rom[185][55] = 16'h002C;
        rom[185][56] = 16'h0004;
        rom[185][57] = 16'h0035;
        rom[185][58] = 16'hFFE4;
        rom[185][59] = 16'hFFED;
        rom[185][60] = 16'h0002;
        rom[185][61] = 16'hFFE1;
        rom[185][62] = 16'hFFBB;
        rom[185][63] = 16'hFFFE;
        rom[185][64] = 16'h0003;
        rom[185][65] = 16'hFFE6;
        rom[185][66] = 16'hFFF8;
        rom[185][67] = 16'hFFDF;
        rom[185][68] = 16'hFFEF;
        rom[185][69] = 16'h001D;
        rom[185][70] = 16'h000B;
        rom[185][71] = 16'h000D;
        rom[185][72] = 16'h000C;
        rom[185][73] = 16'hFFB5;
        rom[185][74] = 16'hFFE7;
        rom[185][75] = 16'h0024;
        rom[185][76] = 16'h0019;
        rom[185][77] = 16'hFFB3;
        rom[185][78] = 16'hFFF4;
        rom[185][79] = 16'hFFBF;
        rom[185][80] = 16'hFFDC;
        rom[185][81] = 16'hFFDB;
        rom[185][82] = 16'hFFE4;
        rom[185][83] = 16'hFFD4;
        rom[185][84] = 16'hFFDC;
        rom[185][85] = 16'hFFCD;
        rom[185][86] = 16'hFFF6;
        rom[185][87] = 16'h000C;
        rom[185][88] = 16'hFFAF;
        rom[185][89] = 16'hFFEF;
        rom[185][90] = 16'hFFF9;
        rom[185][91] = 16'hFFF0;
        rom[185][92] = 16'hFFFC;
        rom[185][93] = 16'hFFDF;
        rom[185][94] = 16'hFFE7;
        rom[185][95] = 16'hFFE8;
        rom[185][96] = 16'h0012;
        rom[185][97] = 16'hFFFF;
        rom[185][98] = 16'hFFFC;
        rom[185][99] = 16'h0006;
        rom[185][100] = 16'h0014;
        rom[185][101] = 16'h0024;
        rom[185][102] = 16'h0037;
        rom[185][103] = 16'h0030;
        rom[185][104] = 16'hFFED;
        rom[185][105] = 16'h0008;
        rom[185][106] = 16'hFFFE;
        rom[185][107] = 16'hFFEC;
        rom[185][108] = 16'hFFE5;
        rom[185][109] = 16'hFFED;
        rom[185][110] = 16'hFFC8;
        rom[185][111] = 16'hFFDF;
        rom[185][112] = 16'h0000;
        rom[185][113] = 16'hFFCC;
        rom[185][114] = 16'h0028;
        rom[185][115] = 16'h000F;
        rom[185][116] = 16'h0013;
        rom[185][117] = 16'hFFFE;
        rom[185][118] = 16'hFFFC;
        rom[185][119] = 16'hFFF5;
        rom[185][120] = 16'hFFEA;
        rom[185][121] = 16'h0017;
        rom[185][122] = 16'hFFFA;
        rom[185][123] = 16'hFFD4;
        rom[185][124] = 16'hFFCB;
        rom[185][125] = 16'hFFC2;
        rom[185][126] = 16'hFFF0;
        rom[185][127] = 16'h001A;
        rom[186][0] = 16'h0016;
        rom[186][1] = 16'hFFD5;
        rom[186][2] = 16'hFFC1;
        rom[186][3] = 16'h000C;
        rom[186][4] = 16'hFFF4;
        rom[186][5] = 16'hFFDF;
        rom[186][6] = 16'h001E;
        rom[186][7] = 16'h0009;
        rom[186][8] = 16'hFFC3;
        rom[186][9] = 16'hFFC6;
        rom[186][10] = 16'hFFD3;
        rom[186][11] = 16'hFFDA;
        rom[186][12] = 16'h001B;
        rom[186][13] = 16'h0029;
        rom[186][14] = 16'hFFEF;
        rom[186][15] = 16'hFFD4;
        rom[186][16] = 16'hFFF1;
        rom[186][17] = 16'h000C;
        rom[186][18] = 16'hFFF7;
        rom[186][19] = 16'hFFF3;
        rom[186][20] = 16'h0010;
        rom[186][21] = 16'hFFE9;
        rom[186][22] = 16'h002A;
        rom[186][23] = 16'hFFC5;
        rom[186][24] = 16'hFFFC;
        rom[186][25] = 16'hFFF1;
        rom[186][26] = 16'h0004;
        rom[186][27] = 16'hFFFE;
        rom[186][28] = 16'h0017;
        rom[186][29] = 16'hFFF0;
        rom[186][30] = 16'h0017;
        rom[186][31] = 16'hFFE6;
        rom[186][32] = 16'hFFCB;
        rom[186][33] = 16'hFFAD;
        rom[186][34] = 16'h0033;
        rom[186][35] = 16'h0010;
        rom[186][36] = 16'h0024;
        rom[186][37] = 16'h0024;
        rom[186][38] = 16'hFFDA;
        rom[186][39] = 16'h0004;
        rom[186][40] = 16'h0027;
        rom[186][41] = 16'hFFD2;
        rom[186][42] = 16'h000C;
        rom[186][43] = 16'hFFF4;
        rom[186][44] = 16'h0002;
        rom[186][45] = 16'hFFC8;
        rom[186][46] = 16'hFFDD;
        rom[186][47] = 16'hFFDE;
        rom[186][48] = 16'h0009;
        rom[186][49] = 16'hFFE5;
        rom[186][50] = 16'hFFD7;
        rom[186][51] = 16'h0026;
        rom[186][52] = 16'hFFD3;
        rom[186][53] = 16'hFFEB;
        rom[186][54] = 16'hFFD0;
        rom[186][55] = 16'hFFFE;
        rom[186][56] = 16'hFFFE;
        rom[186][57] = 16'hFFE0;
        rom[186][58] = 16'hFFED;
        rom[186][59] = 16'hFFF6;
        rom[186][60] = 16'h0013;
        rom[186][61] = 16'hFFEF;
        rom[186][62] = 16'hFFFE;
        rom[186][63] = 16'h0007;
        rom[186][64] = 16'h0024;
        rom[186][65] = 16'h002F;
        rom[186][66] = 16'hFFE8;
        rom[186][67] = 16'hFFFE;
        rom[186][68] = 16'h0026;
        rom[186][69] = 16'h0004;
        rom[186][70] = 16'hFFEA;
        rom[186][71] = 16'hFFF7;
        rom[186][72] = 16'hFFE5;
        rom[186][73] = 16'h0011;
        rom[186][74] = 16'h0011;
        rom[186][75] = 16'hFFC5;
        rom[186][76] = 16'hFFC7;
        rom[186][77] = 16'hFFF3;
        rom[186][78] = 16'hFFFE;
        rom[186][79] = 16'h0006;
        rom[186][80] = 16'h001F;
        rom[186][81] = 16'hFFF5;
        rom[186][82] = 16'hFFC9;
        rom[186][83] = 16'hFFE5;
        rom[186][84] = 16'hFFDE;
        rom[186][85] = 16'hFFE0;
        rom[186][86] = 16'h0009;
        rom[186][87] = 16'hFFFD;
        rom[186][88] = 16'hFFF4;
        rom[186][89] = 16'hFFE7;
        rom[186][90] = 16'hFFF2;
        rom[186][91] = 16'h001B;
        rom[186][92] = 16'h002B;
        rom[186][93] = 16'h000D;
        rom[186][94] = 16'h0003;
        rom[186][95] = 16'h0005;
        rom[186][96] = 16'h0018;
        rom[186][97] = 16'hFFF4;
        rom[186][98] = 16'hFFFE;
        rom[186][99] = 16'h0012;
        rom[186][100] = 16'h0015;
        rom[186][101] = 16'h000A;
        rom[186][102] = 16'h0009;
        rom[186][103] = 16'h000A;
        rom[186][104] = 16'h0035;
        rom[186][105] = 16'hFFC8;
        rom[186][106] = 16'h000A;
        rom[186][107] = 16'hFFBC;
        rom[186][108] = 16'hFFEA;
        rom[186][109] = 16'h0026;
        rom[186][110] = 16'h0007;
        rom[186][111] = 16'hFFF2;
        rom[186][112] = 16'hFFEE;
        rom[186][113] = 16'hFFEA;
        rom[186][114] = 16'hFFF8;
        rom[186][115] = 16'h001A;
        rom[186][116] = 16'hFFC4;
        rom[186][117] = 16'h0001;
        rom[186][118] = 16'hFFD8;
        rom[186][119] = 16'hFFAA;
        rom[186][120] = 16'h0015;
        rom[186][121] = 16'hFFE6;
        rom[186][122] = 16'hFFCC;
        rom[186][123] = 16'hFFF4;
        rom[186][124] = 16'hFFE6;
        rom[186][125] = 16'h001F;
        rom[186][126] = 16'h0008;
        rom[186][127] = 16'h000A;
        rom[187][0] = 16'h0011;
        rom[187][1] = 16'hFFE6;
        rom[187][2] = 16'h000D;
        rom[187][3] = 16'h0019;
        rom[187][4] = 16'hFFCF;
        rom[187][5] = 16'hFFB9;
        rom[187][6] = 16'h0004;
        rom[187][7] = 16'h0009;
        rom[187][8] = 16'hFFCC;
        rom[187][9] = 16'hFFFE;
        rom[187][10] = 16'hFFE3;
        rom[187][11] = 16'hFFEC;
        rom[187][12] = 16'hFFC4;
        rom[187][13] = 16'h0007;
        rom[187][14] = 16'hFFCD;
        rom[187][15] = 16'h0002;
        rom[187][16] = 16'hFFDE;
        rom[187][17] = 16'hFFF3;
        rom[187][18] = 16'h0012;
        rom[187][19] = 16'h0016;
        rom[187][20] = 16'hFFDC;
        rom[187][21] = 16'hFFFD;
        rom[187][22] = 16'hFFE8;
        rom[187][23] = 16'h000F;
        rom[187][24] = 16'h000E;
        rom[187][25] = 16'hFFEA;
        rom[187][26] = 16'hFFF1;
        rom[187][27] = 16'hFFDD;
        rom[187][28] = 16'hFFFE;
        rom[187][29] = 16'hFFFE;
        rom[187][30] = 16'h000E;
        rom[187][31] = 16'h001B;
        rom[187][32] = 16'hFFE2;
        rom[187][33] = 16'h002A;
        rom[187][34] = 16'hFFFA;
        rom[187][35] = 16'hFFEA;
        rom[187][36] = 16'h0001;
        rom[187][37] = 16'hFFDC;
        rom[187][38] = 16'hFFED;
        rom[187][39] = 16'h0033;
        rom[187][40] = 16'hFFEB;
        rom[187][41] = 16'h0011;
        rom[187][42] = 16'hFFE3;
        rom[187][43] = 16'hFFEF;
        rom[187][44] = 16'h0012;
        rom[187][45] = 16'hFFF9;
        rom[187][46] = 16'h0015;
        rom[187][47] = 16'h0032;
        rom[187][48] = 16'hFFC5;
        rom[187][49] = 16'hFFDE;
        rom[187][50] = 16'hFFDA;
        rom[187][51] = 16'h0007;
        rom[187][52] = 16'hFFD8;
        rom[187][53] = 16'hFFD1;
        rom[187][54] = 16'h002B;
        rom[187][55] = 16'hFFD2;
        rom[187][56] = 16'hFFE0;
        rom[187][57] = 16'hFFF2;
        rom[187][58] = 16'h0017;
        rom[187][59] = 16'hFFED;
        rom[187][60] = 16'hFFF7;
        rom[187][61] = 16'h0020;
        rom[187][62] = 16'h0000;
        rom[187][63] = 16'hFFE7;
        rom[187][64] = 16'h001D;
        rom[187][65] = 16'hFFFE;
        rom[187][66] = 16'hFFC8;
        rom[187][67] = 16'hFFCE;
        rom[187][68] = 16'h0002;
        rom[187][69] = 16'hFFDE;
        rom[187][70] = 16'hFFF7;
        rom[187][71] = 16'hFFFD;
        rom[187][72] = 16'h0004;
        rom[187][73] = 16'hFFE5;
        rom[187][74] = 16'h0011;
        rom[187][75] = 16'h001D;
        rom[187][76] = 16'h0000;
        rom[187][77] = 16'hFFDF;
        rom[187][78] = 16'h0017;
        rom[187][79] = 16'hFFF1;
        rom[187][80] = 16'hFFF9;
        rom[187][81] = 16'h001D;
        rom[187][82] = 16'hFFD8;
        rom[187][83] = 16'hFFE8;
        rom[187][84] = 16'hFFD6;
        rom[187][85] = 16'hFFEA;
        rom[187][86] = 16'h002C;
        rom[187][87] = 16'hFFDB;
        rom[187][88] = 16'h0005;
        rom[187][89] = 16'hFFEE;
        rom[187][90] = 16'hFFFB;
        rom[187][91] = 16'hFFF1;
        rom[187][92] = 16'h0003;
        rom[187][93] = 16'h0001;
        rom[187][94] = 16'h001B;
        rom[187][95] = 16'hFFE2;
        rom[187][96] = 16'hFFF4;
        rom[187][97] = 16'hFFF8;
        rom[187][98] = 16'h002F;
        rom[187][99] = 16'h0007;
        rom[187][100] = 16'h0021;
        rom[187][101] = 16'h000F;
        rom[187][102] = 16'hFFE3;
        rom[187][103] = 16'hFFE5;
        rom[187][104] = 16'h001F;
        rom[187][105] = 16'hFFD1;
        rom[187][106] = 16'h0001;
        rom[187][107] = 16'hFFCA;
        rom[187][108] = 16'hFFEF;
        rom[187][109] = 16'h0015;
        rom[187][110] = 16'hFFCF;
        rom[187][111] = 16'hFFFF;
        rom[187][112] = 16'h0010;
        rom[187][113] = 16'hFFE4;
        rom[187][114] = 16'hFFF4;
        rom[187][115] = 16'hFFDB;
        rom[187][116] = 16'hFFDC;
        rom[187][117] = 16'hFFE8;
        rom[187][118] = 16'hFFE1;
        rom[187][119] = 16'h0001;
        rom[187][120] = 16'h0002;
        rom[187][121] = 16'hFFFF;
        rom[187][122] = 16'hFFE1;
        rom[187][123] = 16'hFFF6;
        rom[187][124] = 16'h000C;
        rom[187][125] = 16'h001A;
        rom[187][126] = 16'hFFCD;
        rom[187][127] = 16'hFFB3;
        rom[188][0] = 16'h0014;
        rom[188][1] = 16'hFFF5;
        rom[188][2] = 16'hFFFB;
        rom[188][3] = 16'h0007;
        rom[188][4] = 16'h0005;
        rom[188][5] = 16'h0015;
        rom[188][6] = 16'hFFE1;
        rom[188][7] = 16'hFFD7;
        rom[188][8] = 16'h000F;
        rom[188][9] = 16'hFFFE;
        rom[188][10] = 16'hFFDF;
        rom[188][11] = 16'hFFE5;
        rom[188][12] = 16'hFFE3;
        rom[188][13] = 16'hFFF3;
        rom[188][14] = 16'hFFF7;
        rom[188][15] = 16'h001F;
        rom[188][16] = 16'hFFD5;
        rom[188][17] = 16'hFF97;
        rom[188][18] = 16'hFFFE;
        rom[188][19] = 16'hFFEA;
        rom[188][20] = 16'hFFF4;
        rom[188][21] = 16'h0021;
        rom[188][22] = 16'hFFC9;
        rom[188][23] = 16'hFFE5;
        rom[188][24] = 16'hFFFE;
        rom[188][25] = 16'h0017;
        rom[188][26] = 16'hFFC8;
        rom[188][27] = 16'h0020;
        rom[188][28] = 16'h000E;
        rom[188][29] = 16'h0008;
        rom[188][30] = 16'h0010;
        rom[188][31] = 16'h0001;
        rom[188][32] = 16'hFFEA;
        rom[188][33] = 16'hFFD7;
        rom[188][34] = 16'h0006;
        rom[188][35] = 16'h0014;
        rom[188][36] = 16'hFFCD;
        rom[188][37] = 16'hFFBC;
        rom[188][38] = 16'h000A;
        rom[188][39] = 16'hFFF2;
        rom[188][40] = 16'hFFE1;
        rom[188][41] = 16'h0002;
        rom[188][42] = 16'hFFDA;
        rom[188][43] = 16'h0012;
        rom[188][44] = 16'hFFF4;
        rom[188][45] = 16'hFFD8;
        rom[188][46] = 16'hFFD4;
        rom[188][47] = 16'h000B;
        rom[188][48] = 16'hFFDC;
        rom[188][49] = 16'hFFED;
        rom[188][50] = 16'hFFFC;
        rom[188][51] = 16'h000C;
        rom[188][52] = 16'h0011;
        rom[188][53] = 16'hFFEA;
        rom[188][54] = 16'hFFEC;
        rom[188][55] = 16'h0026;
        rom[188][56] = 16'h000E;
        rom[188][57] = 16'h0000;
        rom[188][58] = 16'hFFE5;
        rom[188][59] = 16'hFFF9;
        rom[188][60] = 16'hFFE0;
        rom[188][61] = 16'h0001;
        rom[188][62] = 16'h0031;
        rom[188][63] = 16'hFFEA;
        rom[188][64] = 16'h0011;
        rom[188][65] = 16'hFFBC;
        rom[188][66] = 16'hFFF1;
        rom[188][67] = 16'h0013;
        rom[188][68] = 16'hFFFD;
        rom[188][69] = 16'h0023;
        rom[188][70] = 16'h0002;
        rom[188][71] = 16'hFFF2;
        rom[188][72] = 16'h0011;
        rom[188][73] = 16'h0025;
        rom[188][74] = 16'hFFE3;
        rom[188][75] = 16'h0027;
        rom[188][76] = 16'hFFD7;
        rom[188][77] = 16'hFFF1;
        rom[188][78] = 16'h0001;
        rom[188][79] = 16'hFFEA;
        rom[188][80] = 16'hFFD0;
        rom[188][81] = 16'hFFC7;
        rom[188][82] = 16'hFFEF;
        rom[188][83] = 16'h001A;
        rom[188][84] = 16'hFFB1;
        rom[188][85] = 16'h0020;
        rom[188][86] = 16'h000B;
        rom[188][87] = 16'hFFE8;
        rom[188][88] = 16'hFFFD;
        rom[188][89] = 16'h0003;
        rom[188][90] = 16'hFFF6;
        rom[188][91] = 16'hFFE9;
        rom[188][92] = 16'hFFE1;
        rom[188][93] = 16'h0007;
        rom[188][94] = 16'hFFE1;
        rom[188][95] = 16'hFFDB;
        rom[188][96] = 16'hFFF0;
        rom[188][97] = 16'hFFB2;
        rom[188][98] = 16'h0020;
        rom[188][99] = 16'hFFBC;
        rom[188][100] = 16'h000B;
        rom[188][101] = 16'hFFFC;
        rom[188][102] = 16'hFFC4;
        rom[188][103] = 16'h0005;
        rom[188][104] = 16'h0014;
        rom[188][105] = 16'hFFE9;
        rom[188][106] = 16'hFFE1;
        rom[188][107] = 16'h0002;
        rom[188][108] = 16'h0002;
        rom[188][109] = 16'hFFFE;
        rom[188][110] = 16'h0018;
        rom[188][111] = 16'h0030;
        rom[188][112] = 16'h000F;
        rom[188][113] = 16'h0032;
        rom[188][114] = 16'hFFFE;
        rom[188][115] = 16'hFFFF;
        rom[188][116] = 16'hFFE3;
        rom[188][117] = 16'hFFE1;
        rom[188][118] = 16'h0024;
        rom[188][119] = 16'hFFDC;
        rom[188][120] = 16'h0010;
        rom[188][121] = 16'h0031;
        rom[188][122] = 16'h000B;
        rom[188][123] = 16'hFFE0;
        rom[188][124] = 16'hFFDA;
        rom[188][125] = 16'h0016;
        rom[188][126] = 16'hFFF9;
        rom[188][127] = 16'hFFFF;
        rom[189][0] = 16'hFFEF;
        rom[189][1] = 16'h001E;
        rom[189][2] = 16'h0001;
        rom[189][3] = 16'h001E;
        rom[189][4] = 16'hFFD1;
        rom[189][5] = 16'hFFE6;
        rom[189][6] = 16'h0020;
        rom[189][7] = 16'hFFF4;
        rom[189][8] = 16'h0002;
        rom[189][9] = 16'hFFC3;
        rom[189][10] = 16'hFFFC;
        rom[189][11] = 16'h0028;
        rom[189][12] = 16'h0041;
        rom[189][13] = 16'hFFE9;
        rom[189][14] = 16'hFFD6;
        rom[189][15] = 16'hFFC9;
        rom[189][16] = 16'h0021;
        rom[189][17] = 16'hFFE4;
        rom[189][18] = 16'h0016;
        rom[189][19] = 16'h0006;
        rom[189][20] = 16'h0016;
        rom[189][21] = 16'hFFE1;
        rom[189][22] = 16'hFFFA;
        rom[189][23] = 16'h0027;
        rom[189][24] = 16'h001A;
        rom[189][25] = 16'hFFD9;
        rom[189][26] = 16'h003A;
        rom[189][27] = 16'hFFD8;
        rom[189][28] = 16'hFFE0;
        rom[189][29] = 16'hFFD4;
        rom[189][30] = 16'hFFDA;
        rom[189][31] = 16'hFFE4;
        rom[189][32] = 16'h0011;
        rom[189][33] = 16'hFFD6;
        rom[189][34] = 16'hFFD7;
        rom[189][35] = 16'hFFD4;
        rom[189][36] = 16'h0008;
        rom[189][37] = 16'hFFEC;
        rom[189][38] = 16'hFFC0;
        rom[189][39] = 16'h000D;
        rom[189][40] = 16'hFFD2;
        rom[189][41] = 16'hFFC5;
        rom[189][42] = 16'h0021;
        rom[189][43] = 16'hFFEA;
        rom[189][44] = 16'h000D;
        rom[189][45] = 16'hFFEF;
        rom[189][46] = 16'h001F;
        rom[189][47] = 16'hFFE5;
        rom[189][48] = 16'h0000;
        rom[189][49] = 16'h001F;
        rom[189][50] = 16'hFFFC;
        rom[189][51] = 16'hFFFE;
        rom[189][52] = 16'hFFEF;
        rom[189][53] = 16'hFFDE;
        rom[189][54] = 16'hFFDC;
        rom[189][55] = 16'hFFC0;
        rom[189][56] = 16'hFFE6;
        rom[189][57] = 16'h003A;
        rom[189][58] = 16'h0016;
        rom[189][59] = 16'h003E;
        rom[189][60] = 16'hFFF5;
        rom[189][61] = 16'hFFFF;
        rom[189][62] = 16'hFFFE;
        rom[189][63] = 16'h0014;
        rom[189][64] = 16'h0002;
        rom[189][65] = 16'hFFFE;
        rom[189][66] = 16'hFFD8;
        rom[189][67] = 16'hFFEA;
        rom[189][68] = 16'hFFD4;
        rom[189][69] = 16'h0019;
        rom[189][70] = 16'hFFC8;
        rom[189][71] = 16'h0009;
        rom[189][72] = 16'h0022;
        rom[189][73] = 16'hFFCF;
        rom[189][74] = 16'hFFF5;
        rom[189][75] = 16'h0006;
        rom[189][76] = 16'h000C;
        rom[189][77] = 16'h0002;
        rom[189][78] = 16'hFFDB;
        rom[189][79] = 16'h001F;
        rom[189][80] = 16'h0045;
        rom[189][81] = 16'h0003;
        rom[189][82] = 16'h0020;
        rom[189][83] = 16'hFFE5;
        rom[189][84] = 16'h0002;
        rom[189][85] = 16'h000A;
        rom[189][86] = 16'h0005;
        rom[189][87] = 16'h0007;
        rom[189][88] = 16'h001B;
        rom[189][89] = 16'hFFB7;
        rom[189][90] = 16'h0032;
        rom[189][91] = 16'h0009;
        rom[189][92] = 16'hFFF4;
        rom[189][93] = 16'h0002;
        rom[189][94] = 16'hFFEE;
        rom[189][95] = 16'hFFE1;
        rom[189][96] = 16'h0002;
        rom[189][97] = 16'h0024;
        rom[189][98] = 16'h0044;
        rom[189][99] = 16'h000C;
        rom[189][100] = 16'hFFFB;
        rom[189][101] = 16'hFFCD;
        rom[189][102] = 16'h000C;
        rom[189][103] = 16'h0023;
        rom[189][104] = 16'hFFF6;
        rom[189][105] = 16'hFFE9;
        rom[189][106] = 16'hFFC4;
        rom[189][107] = 16'hFFEB;
        rom[189][108] = 16'h0012;
        rom[189][109] = 16'hFFD8;
        rom[189][110] = 16'hFFEF;
        rom[189][111] = 16'h0002;
        rom[189][112] = 16'h0001;
        rom[189][113] = 16'h0024;
        rom[189][114] = 16'h0038;
        rom[189][115] = 16'hFFEE;
        rom[189][116] = 16'h000E;
        rom[189][117] = 16'h002E;
        rom[189][118] = 16'h001F;
        rom[189][119] = 16'hFFEF;
        rom[189][120] = 16'h0014;
        rom[189][121] = 16'h0033;
        rom[189][122] = 16'h004B;
        rom[189][123] = 16'hFFD8;
        rom[189][124] = 16'h0001;
        rom[189][125] = 16'h0003;
        rom[189][126] = 16'hFFEA;
        rom[189][127] = 16'h0005;
        rom[190][0] = 16'h0010;
        rom[190][1] = 16'h0033;
        rom[190][2] = 16'hFFCC;
        rom[190][3] = 16'hFFE5;
        rom[190][4] = 16'hFFFB;
        rom[190][5] = 16'h0010;
        rom[190][6] = 16'hFFE8;
        rom[190][7] = 16'h0018;
        rom[190][8] = 16'h0030;
        rom[190][9] = 16'h0015;
        rom[190][10] = 16'h0002;
        rom[190][11] = 16'hFFC1;
        rom[190][12] = 16'h0006;
        rom[190][13] = 16'h0024;
        rom[190][14] = 16'h0027;
        rom[190][15] = 16'hFFE0;
        rom[190][16] = 16'hFFF6;
        rom[190][17] = 16'h0001;
        rom[190][18] = 16'h0009;
        rom[190][19] = 16'hFFE2;
        rom[190][20] = 16'hFFCD;
        rom[190][21] = 16'hFFFE;
        rom[190][22] = 16'hFFEA;
        rom[190][23] = 16'h000B;
        rom[190][24] = 16'h0002;
        rom[190][25] = 16'h0002;
        rom[190][26] = 16'h000C;
        rom[190][27] = 16'hFF9F;
        rom[190][28] = 16'hFFF1;
        rom[190][29] = 16'hFFD2;
        rom[190][30] = 16'h0017;
        rom[190][31] = 16'h0016;
        rom[190][32] = 16'hFFCB;
        rom[190][33] = 16'h001E;
        rom[190][34] = 16'hFFC4;
        rom[190][35] = 16'hFFD8;
        rom[190][36] = 16'h0035;
        rom[190][37] = 16'h000A;
        rom[190][38] = 16'h002E;
        rom[190][39] = 16'hFFA3;
        rom[190][40] = 16'h000B;
        rom[190][41] = 16'hFFEF;
        rom[190][42] = 16'h0002;
        rom[190][43] = 16'h0015;
        rom[190][44] = 16'hFFFC;
        rom[190][45] = 16'hFFC3;
        rom[190][46] = 16'h0022;
        rom[190][47] = 16'h0007;
        rom[190][48] = 16'h0006;
        rom[190][49] = 16'hFFF4;
        rom[190][50] = 16'hFFEC;
        rom[190][51] = 16'h0001;
        rom[190][52] = 16'hFFD7;
        rom[190][53] = 16'h0024;
        rom[190][54] = 16'hFFDE;
        rom[190][55] = 16'hFFF9;
        rom[190][56] = 16'hFFF7;
        rom[190][57] = 16'h001B;
        rom[190][58] = 16'h0031;
        rom[190][59] = 16'h0007;
        rom[190][60] = 16'hFFF0;
        rom[190][61] = 16'hFFED;
        rom[190][62] = 16'hFFDC;
        rom[190][63] = 16'h0041;
        rom[190][64] = 16'hFFF7;
        rom[190][65] = 16'h002E;
        rom[190][66] = 16'h0009;
        rom[190][67] = 16'h0014;
        rom[190][68] = 16'h0013;
        rom[190][69] = 16'hFFE5;
        rom[190][70] = 16'hFFF8;
        rom[190][71] = 16'hFFC1;
        rom[190][72] = 16'hFFF4;
        rom[190][73] = 16'hFFE0;
        rom[190][74] = 16'h0018;
        rom[190][75] = 16'h0029;
        rom[190][76] = 16'hFFE0;
        rom[190][77] = 16'h0030;
        rom[190][78] = 16'hFFD6;
        rom[190][79] = 16'hFFEA;
        rom[190][80] = 16'h0030;
        rom[190][81] = 16'hFFDF;
        rom[190][82] = 16'h0010;
        rom[190][83] = 16'hFFF9;
        rom[190][84] = 16'h0000;
        rom[190][85] = 16'h0011;
        rom[190][86] = 16'hFFFB;
        rom[190][87] = 16'hFFD5;
        rom[190][88] = 16'hFFE1;
        rom[190][89] = 16'hFFF6;
        rom[190][90] = 16'h0021;
        rom[190][91] = 16'hFFE1;
        rom[190][92] = 16'hFFD6;
        rom[190][93] = 16'hFFD2;
        rom[190][94] = 16'hFFEF;
        rom[190][95] = 16'hFFE5;
        rom[190][96] = 16'hFFD7;
        rom[190][97] = 16'hFFD2;
        rom[190][98] = 16'h001E;
        rom[190][99] = 16'h0011;
        rom[190][100] = 16'hFFD4;
        rom[190][101] = 16'hFFF7;
        rom[190][102] = 16'h0024;
        rom[190][103] = 16'hFFE0;
        rom[190][104] = 16'h0006;
        rom[190][105] = 16'h002A;
        rom[190][106] = 16'hFFF9;
        rom[190][107] = 16'hFFC8;
        rom[190][108] = 16'hFFB0;
        rom[190][109] = 16'hFFCB;
        rom[190][110] = 16'hFFD7;
        rom[190][111] = 16'hFFF5;
        rom[190][112] = 16'hFFDF;
        rom[190][113] = 16'h001F;
        rom[190][114] = 16'hFFCA;
        rom[190][115] = 16'hFFCF;
        rom[190][116] = 16'h0000;
        rom[190][117] = 16'h0014;
        rom[190][118] = 16'h0019;
        rom[190][119] = 16'hFFE1;
        rom[190][120] = 16'hFFCE;
        rom[190][121] = 16'hFFFD;
        rom[190][122] = 16'hFFD7;
        rom[190][123] = 16'hFFF4;
        rom[190][124] = 16'hFFF7;
        rom[190][125] = 16'h000C;
        rom[190][126] = 16'hFFF9;
        rom[190][127] = 16'h001F;
        rom[191][0] = 16'hFFF0;
        rom[191][1] = 16'hFFFC;
        rom[191][2] = 16'hFFE7;
        rom[191][3] = 16'hFFBB;
        rom[191][4] = 16'hFFFF;
        rom[191][5] = 16'h0007;
        rom[191][6] = 16'hFFE1;
        rom[191][7] = 16'h001F;
        rom[191][8] = 16'hFFD6;
        rom[191][9] = 16'h0004;
        rom[191][10] = 16'h000B;
        rom[191][11] = 16'h0000;
        rom[191][12] = 16'h000C;
        rom[191][13] = 16'hFFE5;
        rom[191][14] = 16'hFFD2;
        rom[191][15] = 16'h0001;
        rom[191][16] = 16'hFFF9;
        rom[191][17] = 16'h0024;
        rom[191][18] = 16'h0004;
        rom[191][19] = 16'hFFD8;
        rom[191][20] = 16'hFFFC;
        rom[191][21] = 16'h000B;
        rom[191][22] = 16'hFFD8;
        rom[191][23] = 16'hFFEF;
        rom[191][24] = 16'hFFFD;
        rom[191][25] = 16'hFFBF;
        rom[191][26] = 16'hFFE8;
        rom[191][27] = 16'hFFED;
        rom[191][28] = 16'h0004;
        rom[191][29] = 16'h0013;
        rom[191][30] = 16'h001D;
        rom[191][31] = 16'h001B;
        rom[191][32] = 16'h0002;
        rom[191][33] = 16'h0028;
        rom[191][34] = 16'hFFEA;
        rom[191][35] = 16'h0007;
        rom[191][36] = 16'h000C;
        rom[191][37] = 16'hFFFE;
        rom[191][38] = 16'hFFE5;
        rom[191][39] = 16'h002C;
        rom[191][40] = 16'hFFDB;
        rom[191][41] = 16'hFFFC;
        rom[191][42] = 16'hFFF4;
        rom[191][43] = 16'h0029;
        rom[191][44] = 16'h0026;
        rom[191][45] = 16'h0016;
        rom[191][46] = 16'h000B;
        rom[191][47] = 16'h0036;
        rom[191][48] = 16'h000D;
        rom[191][49] = 16'h0007;
        rom[191][50] = 16'h0001;
        rom[191][51] = 16'hFFD6;
        rom[191][52] = 16'hFFEB;
        rom[191][53] = 16'hFFD9;
        rom[191][54] = 16'h0019;
        rom[191][55] = 16'h0015;
        rom[191][56] = 16'h001E;
        rom[191][57] = 16'hFFE8;
        rom[191][58] = 16'h0021;
        rom[191][59] = 16'h0011;
        rom[191][60] = 16'h001E;
        rom[191][61] = 16'hFFF4;
        rom[191][62] = 16'h0002;
        rom[191][63] = 16'hFFF0;
        rom[191][64] = 16'hFFE3;
        rom[191][65] = 16'h000C;
        rom[191][66] = 16'h0003;
        rom[191][67] = 16'hFFDF;
        rom[191][68] = 16'hFFEB;
        rom[191][69] = 16'hFFF9;
        rom[191][70] = 16'hFFC2;
        rom[191][71] = 16'hFFF9;
        rom[191][72] = 16'h0017;
        rom[191][73] = 16'hFFEF;
        rom[191][74] = 16'hFFFC;
        rom[191][75] = 16'h0015;
        rom[191][76] = 16'hFFDF;
        rom[191][77] = 16'h003D;
        rom[191][78] = 16'hFFF8;
        rom[191][79] = 16'h000C;
        rom[191][80] = 16'hFFEE;
        rom[191][81] = 16'h002E;
        rom[191][82] = 16'hFFE6;
        rom[191][83] = 16'h0019;
        rom[191][84] = 16'h0002;
        rom[191][85] = 16'hFFFF;
        rom[191][86] = 16'h000F;
        rom[191][87] = 16'hFFE3;
        rom[191][88] = 16'hFFBF;
        rom[191][89] = 16'h0016;
        rom[191][90] = 16'hFFED;
        rom[191][91] = 16'hFFE4;
        rom[191][92] = 16'hFFC4;
        rom[191][93] = 16'h0028;
        rom[191][94] = 16'h0029;
        rom[191][95] = 16'h0006;
        rom[191][96] = 16'hFFF7;
        rom[191][97] = 16'hFFD2;
        rom[191][98] = 16'h002B;
        rom[191][99] = 16'h0036;
        rom[191][100] = 16'h0022;
        rom[191][101] = 16'hFFFC;
        rom[191][102] = 16'hFFF1;
        rom[191][103] = 16'hFFD9;
        rom[191][104] = 16'hFFDE;
        rom[191][105] = 16'hFFC8;
        rom[191][106] = 16'hFFF4;
        rom[191][107] = 16'h001B;
        rom[191][108] = 16'h000F;
        rom[191][109] = 16'h001A;
        rom[191][110] = 16'hFFF7;
        rom[191][111] = 16'h0002;
        rom[191][112] = 16'h000B;
        rom[191][113] = 16'hFFC8;
        rom[191][114] = 16'h0010;
        rom[191][115] = 16'hFFFE;
        rom[191][116] = 16'h0024;
        rom[191][117] = 16'hFFE3;
        rom[191][118] = 16'h000C;
        rom[191][119] = 16'h001C;
        rom[191][120] = 16'hFFEF;
        rom[191][121] = 16'hFFF6;
        rom[191][122] = 16'hFFEB;
        rom[191][123] = 16'hFFFD;
        rom[191][124] = 16'hFFFE;
        rom[191][125] = 16'hFFDF;
        rom[191][126] = 16'hFFDC;
        rom[191][127] = 16'hFFFC;
        rom[192][0] = 16'hFFF6;
        rom[192][1] = 16'h0005;
        rom[192][2] = 16'h0024;
        rom[192][3] = 16'h0010;
        rom[192][4] = 16'h001F;
        rom[192][5] = 16'h0008;
        rom[192][6] = 16'hFFFE;
        rom[192][7] = 16'h0027;
        rom[192][8] = 16'h0012;
        rom[192][9] = 16'h0012;
        rom[192][10] = 16'h001F;
        rom[192][11] = 16'h000C;
        rom[192][12] = 16'hFFB4;
        rom[192][13] = 16'h0003;
        rom[192][14] = 16'h001A;
        rom[192][15] = 16'h0007;
        rom[192][16] = 16'hFFF2;
        rom[192][17] = 16'h0030;
        rom[192][18] = 16'h0014;
        rom[192][19] = 16'h001A;
        rom[192][20] = 16'h0006;
        rom[192][21] = 16'h000C;
        rom[192][22] = 16'h001B;
        rom[192][23] = 16'h0010;
        rom[192][24] = 16'hFFF9;
        rom[192][25] = 16'hFFEB;
        rom[192][26] = 16'hFFFA;
        rom[192][27] = 16'hFFBE;
        rom[192][28] = 16'hFFE5;
        rom[192][29] = 16'h0013;
        rom[192][30] = 16'h0008;
        rom[192][31] = 16'hFFC4;
        rom[192][32] = 16'h0000;
        rom[192][33] = 16'h000C;
        rom[192][34] = 16'h000B;
        rom[192][35] = 16'hFFA0;
        rom[192][36] = 16'hFFFD;
        rom[192][37] = 16'h0002;
        rom[192][38] = 16'h0008;
        rom[192][39] = 16'hFFF4;
        rom[192][40] = 16'h0024;
        rom[192][41] = 16'h0003;
        rom[192][42] = 16'hFFF9;
        rom[192][43] = 16'hFFB1;
        rom[192][44] = 16'hFFC3;
        rom[192][45] = 16'hFFE9;
        rom[192][46] = 16'h0009;
        rom[192][47] = 16'hFFE8;
        rom[192][48] = 16'hFFD9;
        rom[192][49] = 16'hFFF7;
        rom[192][50] = 16'hFFE9;
        rom[192][51] = 16'h0013;
        rom[192][52] = 16'hFFD6;
        rom[192][53] = 16'hFFD4;
        rom[192][54] = 16'hFFD7;
        rom[192][55] = 16'hFFB6;
        rom[192][56] = 16'h0027;
        rom[192][57] = 16'h000A;
        rom[192][58] = 16'hFFD9;
        rom[192][59] = 16'hFFFE;
        rom[192][60] = 16'hFFF3;
        rom[192][61] = 16'hFFFE;
        rom[192][62] = 16'hFFD7;
        rom[192][63] = 16'h002C;
        rom[192][64] = 16'h0016;
        rom[192][65] = 16'hFFF3;
        rom[192][66] = 16'h0017;
        rom[192][67] = 16'hFFFE;
        rom[192][68] = 16'h002A;
        rom[192][69] = 16'hFFF5;
        rom[192][70] = 16'h000C;
        rom[192][71] = 16'hFFEF;
        rom[192][72] = 16'h000F;
        rom[192][73] = 16'h0015;
        rom[192][74] = 16'h001B;
        rom[192][75] = 16'h001C;
        rom[192][76] = 16'h0002;
        rom[192][77] = 16'h0005;
        rom[192][78] = 16'hFFF2;
        rom[192][79] = 16'hFFB9;
        rom[192][80] = 16'h0010;
        rom[192][81] = 16'hFFC6;
        rom[192][82] = 16'hFFFB;
        rom[192][83] = 16'hFFCE;
        rom[192][84] = 16'h000C;
        rom[192][85] = 16'hFFFC;
        rom[192][86] = 16'h0029;
        rom[192][87] = 16'h0013;
        rom[192][88] = 16'h000C;
        rom[192][89] = 16'hFFDC;
        rom[192][90] = 16'h001C;
        rom[192][91] = 16'hFFBF;
        rom[192][92] = 16'hFFFB;
        rom[192][93] = 16'hFFBD;
        rom[192][94] = 16'h0009;
        rom[192][95] = 16'hFFF9;
        rom[192][96] = 16'hFFE3;
        rom[192][97] = 16'h0007;
        rom[192][98] = 16'hFFDE;
        rom[192][99] = 16'hFFB4;
        rom[192][100] = 16'h0021;
        rom[192][101] = 16'hFFE7;
        rom[192][102] = 16'hFFDF;
        rom[192][103] = 16'hFFFD;
        rom[192][104] = 16'hFFF3;
        rom[192][105] = 16'h0008;
        rom[192][106] = 16'h0017;
        rom[192][107] = 16'hFFA6;
        rom[192][108] = 16'hFFF9;
        rom[192][109] = 16'hFFD4;
        rom[192][110] = 16'h000B;
        rom[192][111] = 16'hFFCF;
        rom[192][112] = 16'hFFF4;
        rom[192][113] = 16'h000C;
        rom[192][114] = 16'hFFF4;
        rom[192][115] = 16'hFFE1;
        rom[192][116] = 16'h0009;
        rom[192][117] = 16'hFFFD;
        rom[192][118] = 16'hFFDC;
        rom[192][119] = 16'h0010;
        rom[192][120] = 16'h000D;
        rom[192][121] = 16'h002E;
        rom[192][122] = 16'hFFF4;
        rom[192][123] = 16'hFFF4;
        rom[192][124] = 16'hFFF4;
        rom[192][125] = 16'h0002;
        rom[192][126] = 16'hFFE2;
        rom[192][127] = 16'h0001;
        rom[193][0] = 16'h0011;
        rom[193][1] = 16'hFFF1;
        rom[193][2] = 16'h0007;
        rom[193][3] = 16'hFFEF;
        rom[193][4] = 16'h002D;
        rom[193][5] = 16'h0010;
        rom[193][6] = 16'h0000;
        rom[193][7] = 16'h0019;
        rom[193][8] = 16'h002F;
        rom[193][9] = 16'hFFDE;
        rom[193][10] = 16'hFFEA;
        rom[193][11] = 16'hFFCC;
        rom[193][12] = 16'hFFFB;
        rom[193][13] = 16'hFFF4;
        rom[193][14] = 16'hFFEC;
        rom[193][15] = 16'h0009;
        rom[193][16] = 16'hFFF1;
        rom[193][17] = 16'h001F;
        rom[193][18] = 16'hFFD8;
        rom[193][19] = 16'hFFE0;
        rom[193][20] = 16'hFFDF;
        rom[193][21] = 16'h0001;
        rom[193][22] = 16'h000C;
        rom[193][23] = 16'hFFBB;
        rom[193][24] = 16'hFFEE;
        rom[193][25] = 16'hFFE7;
        rom[193][26] = 16'hFFE1;
        rom[193][27] = 16'hFFEA;
        rom[193][28] = 16'hFFBF;
        rom[193][29] = 16'hFFEE;
        rom[193][30] = 16'h0002;
        rom[193][31] = 16'h001E;
        rom[193][32] = 16'hFFE9;
        rom[193][33] = 16'h0018;
        rom[193][34] = 16'hFFFC;
        rom[193][35] = 16'hFFCF;
        rom[193][36] = 16'hFFCC;
        rom[193][37] = 16'hFFF3;
        rom[193][38] = 16'hFFD7;
        rom[193][39] = 16'hFFF7;
        rom[193][40] = 16'hFFF3;
        rom[193][41] = 16'hFFE0;
        rom[193][42] = 16'hFFF8;
        rom[193][43] = 16'hFFFE;
        rom[193][44] = 16'h0016;
        rom[193][45] = 16'h001B;
        rom[193][46] = 16'hFFB3;
        rom[193][47] = 16'h0015;
        rom[193][48] = 16'hFFE6;
        rom[193][49] = 16'h000E;
        rom[193][50] = 16'h0002;
        rom[193][51] = 16'h0024;
        rom[193][52] = 16'h0020;
        rom[193][53] = 16'h003D;
        rom[193][54] = 16'hFFFA;
        rom[193][55] = 16'hFFE0;
        rom[193][56] = 16'h000A;
        rom[193][57] = 16'h0012;
        rom[193][58] = 16'h0025;
        rom[193][59] = 16'hFFC2;
        rom[193][60] = 16'hFFCD;
        rom[193][61] = 16'hFFF1;
        rom[193][62] = 16'hFFD7;
        rom[193][63] = 16'h000A;
        rom[193][64] = 16'hFFF1;
        rom[193][65] = 16'hFFFF;
        rom[193][66] = 16'h0019;
        rom[193][67] = 16'h0005;
        rom[193][68] = 16'h001B;
        rom[193][69] = 16'h0016;
        rom[193][70] = 16'h0003;
        rom[193][71] = 16'h0011;
        rom[193][72] = 16'h0007;
        rom[193][73] = 16'h000F;
        rom[193][74] = 16'h0016;
        rom[193][75] = 16'hFFDD;
        rom[193][76] = 16'h0003;
        rom[193][77] = 16'hFFF2;
        rom[193][78] = 16'h0001;
        rom[193][79] = 16'hFFEB;
        rom[193][80] = 16'h001A;
        rom[193][81] = 16'h000C;
        rom[193][82] = 16'hFFDB;
        rom[193][83] = 16'hFFF6;
        rom[193][84] = 16'hFFDC;
        rom[193][85] = 16'hFFEC;
        rom[193][86] = 16'hFFD6;
        rom[193][87] = 16'hFFF9;
        rom[193][88] = 16'h0010;
        rom[193][89] = 16'h001D;
        rom[193][90] = 16'hFFE7;
        rom[193][91] = 16'hFFE5;
        rom[193][92] = 16'hFFE7;
        rom[193][93] = 16'hFFE4;
        rom[193][94] = 16'h0011;
        rom[193][95] = 16'hFFE8;
        rom[193][96] = 16'h001F;
        rom[193][97] = 16'h0023;
        rom[193][98] = 16'h000C;
        rom[193][99] = 16'hFFF4;
        rom[193][100] = 16'hFFFF;
        rom[193][101] = 16'hFFD6;
        rom[193][102] = 16'h0011;
        rom[193][103] = 16'h0009;
        rom[193][104] = 16'h0050;
        rom[193][105] = 16'hFFEA;
        rom[193][106] = 16'hFFF4;
        rom[193][107] = 16'h0014;
        rom[193][108] = 16'hFFFD;
        rom[193][109] = 16'hFFE2;
        rom[193][110] = 16'hFFD1;
        rom[193][111] = 16'hFFD6;
        rom[193][112] = 16'hFFE8;
        rom[193][113] = 16'hFFEB;
        rom[193][114] = 16'hFFDC;
        rom[193][115] = 16'hFFFF;
        rom[193][116] = 16'hFFB5;
        rom[193][117] = 16'hFFF8;
        rom[193][118] = 16'hFFF3;
        rom[193][119] = 16'h000C;
        rom[193][120] = 16'hFFFE;
        rom[193][121] = 16'hFFE3;
        rom[193][122] = 16'hFFCF;
        rom[193][123] = 16'hFF9E;
        rom[193][124] = 16'h000D;
        rom[193][125] = 16'h000B;
        rom[193][126] = 16'h0020;
        rom[193][127] = 16'h0015;
        rom[194][0] = 16'h0025;
        rom[194][1] = 16'h0012;
        rom[194][2] = 16'hFFE2;
        rom[194][3] = 16'h001A;
        rom[194][4] = 16'h0005;
        rom[194][5] = 16'hFFE4;
        rom[194][6] = 16'hFFDD;
        rom[194][7] = 16'h001F;
        rom[194][8] = 16'h0007;
        rom[194][9] = 16'h0017;
        rom[194][10] = 16'h0005;
        rom[194][11] = 16'h001E;
        rom[194][12] = 16'hFFFF;
        rom[194][13] = 16'hFFF9;
        rom[194][14] = 16'hFFFA;
        rom[194][15] = 16'h0006;
        rom[194][16] = 16'hFFAC;
        rom[194][17] = 16'h000C;
        rom[194][18] = 16'h000A;
        rom[194][19] = 16'hFFC7;
        rom[194][20] = 16'hFFDF;
        rom[194][21] = 16'hFFF1;
        rom[194][22] = 16'h000D;
        rom[194][23] = 16'h001D;
        rom[194][24] = 16'hFFF2;
        rom[194][25] = 16'hFFDA;
        rom[194][26] = 16'hFFFA;
        rom[194][27] = 16'hFFF8;
        rom[194][28] = 16'h0012;
        rom[194][29] = 16'h0002;
        rom[194][30] = 16'hFFEE;
        rom[194][31] = 16'hFFB9;
        rom[194][32] = 16'h0011;
        rom[194][33] = 16'h001D;
        rom[194][34] = 16'hFFE0;
        rom[194][35] = 16'h0021;
        rom[194][36] = 16'hFFFB;
        rom[194][37] = 16'h0007;
        rom[194][38] = 16'h0014;
        rom[194][39] = 16'h0004;
        rom[194][40] = 16'hFFF2;
        rom[194][41] = 16'h000C;
        rom[194][42] = 16'h0002;
        rom[194][43] = 16'h0008;
        rom[194][44] = 16'hFFD2;
        rom[194][45] = 16'h0017;
        rom[194][46] = 16'hFFF9;
        rom[194][47] = 16'hFFE5;
        rom[194][48] = 16'hFFE4;
        rom[194][49] = 16'h0006;
        rom[194][50] = 16'hFFF2;
        rom[194][51] = 16'hFFEB;
        rom[194][52] = 16'h001B;
        rom[194][53] = 16'h001B;
        rom[194][54] = 16'hFFF7;
        rom[194][55] = 16'hFFFD;
        rom[194][56] = 16'hFFFB;
        rom[194][57] = 16'h0001;
        rom[194][58] = 16'hFFF4;
        rom[194][59] = 16'h0016;
        rom[194][60] = 16'h0064;
        rom[194][61] = 16'hFFDA;
        rom[194][62] = 16'h002F;
        rom[194][63] = 16'hFFEF;
        rom[194][64] = 16'h000F;
        rom[194][65] = 16'h0016;
        rom[194][66] = 16'hFFDA;
        rom[194][67] = 16'h0011;
        rom[194][68] = 16'h0024;
        rom[194][69] = 16'h0016;
        rom[194][70] = 16'hFFF3;
        rom[194][71] = 16'h001A;
        rom[194][72] = 16'hFFDD;
        rom[194][73] = 16'h0016;
        rom[194][74] = 16'hFFEA;
        rom[194][75] = 16'h0005;
        rom[194][76] = 16'hFFEF;
        rom[194][77] = 16'h0003;
        rom[194][78] = 16'hFFC1;
        rom[194][79] = 16'hFFFB;
        rom[194][80] = 16'h0017;
        rom[194][81] = 16'hFFB8;
        rom[194][82] = 16'hFFDF;
        rom[194][83] = 16'h0003;
        rom[194][84] = 16'h0026;
        rom[194][85] = 16'hFFDC;
        rom[194][86] = 16'hFFFB;
        rom[194][87] = 16'hFFEE;
        rom[194][88] = 16'hFFB9;
        rom[194][89] = 16'hFFFF;
        rom[194][90] = 16'hFFD4;
        rom[194][91] = 16'hFFD4;
        rom[194][92] = 16'hFFF6;
        rom[194][93] = 16'h0007;
        rom[194][94] = 16'h000A;
        rom[194][95] = 16'h0016;
        rom[194][96] = 16'h0016;
        rom[194][97] = 16'h001A;
        rom[194][98] = 16'hFFB8;
        rom[194][99] = 16'hFFE5;
        rom[194][100] = 16'h0032;
        rom[194][101] = 16'hFFDB;
        rom[194][102] = 16'h0024;
        rom[194][103] = 16'h000F;
        rom[194][104] = 16'hFFED;
        rom[194][105] = 16'h001B;
        rom[194][106] = 16'hFFDF;
        rom[194][107] = 16'h0030;
        rom[194][108] = 16'h0017;
        rom[194][109] = 16'h0014;
        rom[194][110] = 16'hFFE4;
        rom[194][111] = 16'hFFDA;
        rom[194][112] = 16'hFFF8;
        rom[194][113] = 16'hFFB8;
        rom[194][114] = 16'hFFEC;
        rom[194][115] = 16'hFFFC;
        rom[194][116] = 16'h0008;
        rom[194][117] = 16'h000C;
        rom[194][118] = 16'hFFEB;
        rom[194][119] = 16'hFFF4;
        rom[194][120] = 16'h0000;
        rom[194][121] = 16'hFFF4;
        rom[194][122] = 16'h000A;
        rom[194][123] = 16'hFFEA;
        rom[194][124] = 16'hFFD5;
        rom[194][125] = 16'h0007;
        rom[194][126] = 16'h0042;
        rom[194][127] = 16'h0015;
        rom[195][0] = 16'hFFE9;
        rom[195][1] = 16'hFFEF;
        rom[195][2] = 16'h000A;
        rom[195][3] = 16'hFFFA;
        rom[195][4] = 16'h0019;
        rom[195][5] = 16'h0004;
        rom[195][6] = 16'hFFC4;
        rom[195][7] = 16'hFFC1;
        rom[195][8] = 16'h001A;
        rom[195][9] = 16'hFFF4;
        rom[195][10] = 16'hFFD3;
        rom[195][11] = 16'hFFBD;
        rom[195][12] = 16'hFFF9;
        rom[195][13] = 16'h001B;
        rom[195][14] = 16'hFFEC;
        rom[195][15] = 16'h002C;
        rom[195][16] = 16'h000B;
        rom[195][17] = 16'hFFD2;
        rom[195][18] = 16'hFFBF;
        rom[195][19] = 16'hFFF7;
        rom[195][20] = 16'hFFC2;
        rom[195][21] = 16'h0001;
        rom[195][22] = 16'hFFDC;
        rom[195][23] = 16'hFFD9;
        rom[195][24] = 16'h000E;
        rom[195][25] = 16'hFFDC;
        rom[195][26] = 16'hFFF8;
        rom[195][27] = 16'hFFF5;
        rom[195][28] = 16'h0005;
        rom[195][29] = 16'hFFDE;
        rom[195][30] = 16'h0003;
        rom[195][31] = 16'hFFC5;
        rom[195][32] = 16'h000C;
        rom[195][33] = 16'hFFB4;
        rom[195][34] = 16'hFFE5;
        rom[195][35] = 16'h001E;
        rom[195][36] = 16'hFFC4;
        rom[195][37] = 16'hFFED;
        rom[195][38] = 16'h0000;
        rom[195][39] = 16'h000A;
        rom[195][40] = 16'hFFDC;
        rom[195][41] = 16'h001B;
        rom[195][42] = 16'hFFD8;
        rom[195][43] = 16'h002C;
        rom[195][44] = 16'hFFF3;
        rom[195][45] = 16'h0021;
        rom[195][46] = 16'hFFDC;
        rom[195][47] = 16'hFFF4;
        rom[195][48] = 16'h0004;
        rom[195][49] = 16'h0000;
        rom[195][50] = 16'h000E;
        rom[195][51] = 16'hFFEA;
        rom[195][52] = 16'h0007;
        rom[195][53] = 16'h001B;
        rom[195][54] = 16'h0005;
        rom[195][55] = 16'h0014;
        rom[195][56] = 16'h0004;
        rom[195][57] = 16'hFFFD;
        rom[195][58] = 16'hFFFF;
        rom[195][59] = 16'hFFDC;
        rom[195][60] = 16'h0016;
        rom[195][61] = 16'hFFF9;
        rom[195][62] = 16'h000C;
        rom[195][63] = 16'hFFF2;
        rom[195][64] = 16'h0016;
        rom[195][65] = 16'hFFD3;
        rom[195][66] = 16'h0007;
        rom[195][67] = 16'hFFFC;
        rom[195][68] = 16'hFFE3;
        rom[195][69] = 16'h0027;
        rom[195][70] = 16'h0001;
        rom[195][71] = 16'h0003;
        rom[195][72] = 16'hFFF2;
        rom[195][73] = 16'h0016;
        rom[195][74] = 16'hFFCA;
        rom[195][75] = 16'hFFE3;
        rom[195][76] = 16'h0039;
        rom[195][77] = 16'h000B;
        rom[195][78] = 16'h000E;
        rom[195][79] = 16'hFFE1;
        rom[195][80] = 16'hFFEB;
        rom[195][81] = 16'hFFF3;
        rom[195][82] = 16'hFFE0;
        rom[195][83] = 16'h000A;
        rom[195][84] = 16'h0025;
        rom[195][85] = 16'h000C;
        rom[195][86] = 16'hFFEA;
        rom[195][87] = 16'h0013;
        rom[195][88] = 16'hFFF2;
        rom[195][89] = 16'h0018;
        rom[195][90] = 16'h0003;
        rom[195][91] = 16'hFFF1;
        rom[195][92] = 16'h0007;
        rom[195][93] = 16'hFFC7;
        rom[195][94] = 16'hFFBD;
        rom[195][95] = 16'hFFDB;
        rom[195][96] = 16'h0024;
        rom[195][97] = 16'hFFF5;
        rom[195][98] = 16'hFFF1;
        rom[195][99] = 16'hFFEB;
        rom[195][100] = 16'hFFD7;
        rom[195][101] = 16'h000C;
        rom[195][102] = 16'hFFF0;
        rom[195][103] = 16'hFFF5;
        rom[195][104] = 16'h0008;
        rom[195][105] = 16'hFFC6;
        rom[195][106] = 16'h0009;
        rom[195][107] = 16'h000B;
        rom[195][108] = 16'h0006;
        rom[195][109] = 16'hFFEA;
        rom[195][110] = 16'h0007;
        rom[195][111] = 16'hFFEF;
        rom[195][112] = 16'hFFBD;
        rom[195][113] = 16'h0004;
        rom[195][114] = 16'hFFE5;
        rom[195][115] = 16'hFFD6;
        rom[195][116] = 16'hFFDB;
        rom[195][117] = 16'hFFFE;
        rom[195][118] = 16'h001D;
        rom[195][119] = 16'hFFF9;
        rom[195][120] = 16'h001F;
        rom[195][121] = 16'hFFE0;
        rom[195][122] = 16'h0002;
        rom[195][123] = 16'h000C;
        rom[195][124] = 16'h0003;
        rom[195][125] = 16'h000F;
        rom[195][126] = 16'hFFFD;
        rom[195][127] = 16'h0007;
        rom[196][0] = 16'h0023;
        rom[196][1] = 16'h000C;
        rom[196][2] = 16'h0000;
        rom[196][3] = 16'h0039;
        rom[196][4] = 16'hFFF6;
        rom[196][5] = 16'hFFFF;
        rom[196][6] = 16'h002A;
        rom[196][7] = 16'h0028;
        rom[196][8] = 16'hFFF7;
        rom[196][9] = 16'h0034;
        rom[196][10] = 16'h002B;
        rom[196][11] = 16'hFFCC;
        rom[196][12] = 16'hFFDA;
        rom[196][13] = 16'h000A;
        rom[196][14] = 16'h0003;
        rom[196][15] = 16'hFFEB;
        rom[196][16] = 16'hFFE1;
        rom[196][17] = 16'h0028;
        rom[196][18] = 16'h000D;
        rom[196][19] = 16'h0003;
        rom[196][20] = 16'hFFF2;
        rom[196][21] = 16'hFFE5;
        rom[196][22] = 16'h0024;
        rom[196][23] = 16'h0039;
        rom[196][24] = 16'hFFE7;
        rom[196][25] = 16'h0011;
        rom[196][26] = 16'h0010;
        rom[196][27] = 16'h0006;
        rom[196][28] = 16'hFFFC;
        rom[196][29] = 16'h000A;
        rom[196][30] = 16'hFFFD;
        rom[196][31] = 16'h0016;
        rom[196][32] = 16'h0005;
        rom[196][33] = 16'hFFF7;
        rom[196][34] = 16'h0007;
        rom[196][35] = 16'h0019;
        rom[196][36] = 16'hFFFA;
        rom[196][37] = 16'hFFE4;
        rom[196][38] = 16'h0011;
        rom[196][39] = 16'h0029;
        rom[196][40] = 16'hFFFE;
        rom[196][41] = 16'h000E;
        rom[196][42] = 16'hFFE9;
        rom[196][43] = 16'hFFD4;
        rom[196][44] = 16'h001E;
        rom[196][45] = 16'h002B;
        rom[196][46] = 16'h001B;
        rom[196][47] = 16'h0014;
        rom[196][48] = 16'h002A;
        rom[196][49] = 16'hFFEA;
        rom[196][50] = 16'h002A;
        rom[196][51] = 16'hFFF4;
        rom[196][52] = 16'hFFF5;
        rom[196][53] = 16'h0004;
        rom[196][54] = 16'h000F;
        rom[196][55] = 16'h0019;
        rom[196][56] = 16'hFFD5;
        rom[196][57] = 16'h000C;
        rom[196][58] = 16'hFFE8;
        rom[196][59] = 16'h000B;
        rom[196][60] = 16'hFFEA;
        rom[196][61] = 16'hFFE9;
        rom[196][62] = 16'hFFF3;
        rom[196][63] = 16'h0024;
        rom[196][64] = 16'hFFFC;
        rom[196][65] = 16'h0007;
        rom[196][66] = 16'hFFDB;
        rom[196][67] = 16'hFFBA;
        rom[196][68] = 16'h0017;
        rom[196][69] = 16'hFFE1;
        rom[196][70] = 16'h0023;
        rom[196][71] = 16'hFFDA;
        rom[196][72] = 16'hFFEF;
        rom[196][73] = 16'hFFD5;
        rom[196][74] = 16'h0002;
        rom[196][75] = 16'h0000;
        rom[196][76] = 16'hFFE5;
        rom[196][77] = 16'h000B;
        rom[196][78] = 16'hFFD6;
        rom[196][79] = 16'hFFC4;
        rom[196][80] = 16'hFFF6;
        rom[196][81] = 16'h000A;
        rom[196][82] = 16'hFFED;
        rom[196][83] = 16'h001E;
        rom[196][84] = 16'h0003;
        rom[196][85] = 16'h0038;
        rom[196][86] = 16'h0015;
        rom[196][87] = 16'hFFD1;
        rom[196][88] = 16'h0026;
        rom[196][89] = 16'h0005;
        rom[196][90] = 16'hFFD1;
        rom[196][91] = 16'hFFEA;
        rom[196][92] = 16'hFFDF;
        rom[196][93] = 16'h0007;
        rom[196][94] = 16'hFFF3;
        rom[196][95] = 16'h001C;
        rom[196][96] = 16'hFFFE;
        rom[196][97] = 16'hFFF2;
        rom[196][98] = 16'hFFD0;
        rom[196][99] = 16'h000D;
        rom[196][100] = 16'h000D;
        rom[196][101] = 16'h0004;
        rom[196][102] = 16'hFFDB;
        rom[196][103] = 16'h0004;
        rom[196][104] = 16'hFFC8;
        rom[196][105] = 16'hFFC6;
        rom[196][106] = 16'hFFF8;
        rom[196][107] = 16'hFFC3;
        rom[196][108] = 16'hFFF5;
        rom[196][109] = 16'h001B;
        rom[196][110] = 16'hFFE9;
        rom[196][111] = 16'hFFAB;
        rom[196][112] = 16'hFFF5;
        rom[196][113] = 16'h002E;
        rom[196][114] = 16'hFFC8;
        rom[196][115] = 16'h0043;
        rom[196][116] = 16'h002A;
        rom[196][117] = 16'h000C;
        rom[196][118] = 16'hFFF3;
        rom[196][119] = 16'h001C;
        rom[196][120] = 16'hFFE7;
        rom[196][121] = 16'hFFF9;
        rom[196][122] = 16'hFFC4;
        rom[196][123] = 16'hFFE6;
        rom[196][124] = 16'hFFF1;
        rom[196][125] = 16'hFFE0;
        rom[196][126] = 16'hFFF4;
        rom[196][127] = 16'hFFE0;
        rom[197][0] = 16'h002C;
        rom[197][1] = 16'hFFF9;
        rom[197][2] = 16'hFFE3;
        rom[197][3] = 16'h0032;
        rom[197][4] = 16'hFFE5;
        rom[197][5] = 16'hFFE5;
        rom[197][6] = 16'hFFD8;
        rom[197][7] = 16'h0019;
        rom[197][8] = 16'hFFED;
        rom[197][9] = 16'hFFFA;
        rom[197][10] = 16'hFFEF;
        rom[197][11] = 16'h002E;
        rom[197][12] = 16'h0009;
        rom[197][13] = 16'h0010;
        rom[197][14] = 16'hFFFC;
        rom[197][15] = 16'h001B;
        rom[197][16] = 16'hFFE0;
        rom[197][17] = 16'h0004;
        rom[197][18] = 16'h0018;
        rom[197][19] = 16'hFFE5;
        rom[197][20] = 16'hFFE8;
        rom[197][21] = 16'hFFFB;
        rom[197][22] = 16'h0004;
        rom[197][23] = 16'h001D;
        rom[197][24] = 16'hFFF9;
        rom[197][25] = 16'hFFC1;
        rom[197][26] = 16'hFFBB;
        rom[197][27] = 16'hFFDD;
        rom[197][28] = 16'h0022;
        rom[197][29] = 16'h0001;
        rom[197][30] = 16'hFFF9;
        rom[197][31] = 16'h000A;
        rom[197][32] = 16'h0003;
        rom[197][33] = 16'h0001;
        rom[197][34] = 16'hFFFF;
        rom[197][35] = 16'h0012;
        rom[197][36] = 16'h0017;
        rom[197][37] = 16'h0009;
        rom[197][38] = 16'h001B;
        rom[197][39] = 16'hFFFE;
        rom[197][40] = 16'hFFFC;
        rom[197][41] = 16'hFFF4;
        rom[197][42] = 16'h0007;
        rom[197][43] = 16'h0006;
        rom[197][44] = 16'h000C;
        rom[197][45] = 16'hFFE3;
        rom[197][46] = 16'h002C;
        rom[197][47] = 16'hFFF4;
        rom[197][48] = 16'hFFDB;
        rom[197][49] = 16'hFFCD;
        rom[197][50] = 16'hFFF7;
        rom[197][51] = 16'hFFDC;
        rom[197][52] = 16'hFFD4;
        rom[197][53] = 16'h0004;
        rom[197][54] = 16'h0008;
        rom[197][55] = 16'hFFE9;
        rom[197][56] = 16'hFFCC;
        rom[197][57] = 16'h0016;
        rom[197][58] = 16'hFFD9;
        rom[197][59] = 16'h002D;
        rom[197][60] = 16'hFFF9;
        rom[197][61] = 16'hFFE9;
        rom[197][62] = 16'hFFEE;
        rom[197][63] = 16'hFFE5;
        rom[197][64] = 16'hFFF6;
        rom[197][65] = 16'h0007;
        rom[197][66] = 16'hFFE5;
        rom[197][67] = 16'hFFB8;
        rom[197][68] = 16'h0005;
        rom[197][69] = 16'hFFEB;
        rom[197][70] = 16'h0012;
        rom[197][71] = 16'hFFDE;
        rom[197][72] = 16'h0002;
        rom[197][73] = 16'hFFD2;
        rom[197][74] = 16'h0002;
        rom[197][75] = 16'hFFEC;
        rom[197][76] = 16'h000A;
        rom[197][77] = 16'h0007;
        rom[197][78] = 16'hFFED;
        rom[197][79] = 16'hFFEB;
        rom[197][80] = 16'hFFEE;
        rom[197][81] = 16'hFFFE;
        rom[197][82] = 16'hFFF9;
        rom[197][83] = 16'h0025;
        rom[197][84] = 16'h0017;
        rom[197][85] = 16'h0010;
        rom[197][86] = 16'h0007;
        rom[197][87] = 16'hFFE5;
        rom[197][88] = 16'hFFCA;
        rom[197][89] = 16'h003F;
        rom[197][90] = 16'hFFF9;
        rom[197][91] = 16'hFFD5;
        rom[197][92] = 16'h000E;
        rom[197][93] = 16'h0027;
        rom[197][94] = 16'hFFF0;
        rom[197][95] = 16'h0038;
        rom[197][96] = 16'h0018;
        rom[197][97] = 16'hFFFB;
        rom[197][98] = 16'hFFD2;
        rom[197][99] = 16'h0002;
        rom[197][100] = 16'hFFEF;
        rom[197][101] = 16'hFFDC;
        rom[197][102] = 16'hFFCE;
        rom[197][103] = 16'h0025;
        rom[197][104] = 16'hFFE3;
        rom[197][105] = 16'hFFF4;
        rom[197][106] = 16'h0009;
        rom[197][107] = 16'h0015;
        rom[197][108] = 16'hFFE8;
        rom[197][109] = 16'h0021;
        rom[197][110] = 16'h0029;
        rom[197][111] = 16'hFFE0;
        rom[197][112] = 16'hFFFE;
        rom[197][113] = 16'hFFEC;
        rom[197][114] = 16'hFFEA;
        rom[197][115] = 16'h0013;
        rom[197][116] = 16'h0017;
        rom[197][117] = 16'h0007;
        rom[197][118] = 16'h0010;
        rom[197][119] = 16'hFFEC;
        rom[197][120] = 16'h0024;
        rom[197][121] = 16'h0014;
        rom[197][122] = 16'h000C;
        rom[197][123] = 16'h0015;
        rom[197][124] = 16'h0021;
        rom[197][125] = 16'h0011;
        rom[197][126] = 16'hFFF5;
        rom[197][127] = 16'hFFF6;
        rom[198][0] = 16'hFFE1;
        rom[198][1] = 16'h0006;
        rom[198][2] = 16'h0010;
        rom[198][3] = 16'hFFE6;
        rom[198][4] = 16'h0012;
        rom[198][5] = 16'hFFF1;
        rom[198][6] = 16'h001D;
        rom[198][7] = 16'hFFDC;
        rom[198][8] = 16'h000B;
        rom[198][9] = 16'h001C;
        rom[198][10] = 16'hFFDC;
        rom[198][11] = 16'h0030;
        rom[198][12] = 16'h0007;
        rom[198][13] = 16'hFFF0;
        rom[198][14] = 16'hFFD7;
        rom[198][15] = 16'h0010;
        rom[198][16] = 16'h0003;
        rom[198][17] = 16'hFFC2;
        rom[198][18] = 16'hFFAB;
        rom[198][19] = 16'hFFD8;
        rom[198][20] = 16'h0012;
        rom[198][21] = 16'h0011;
        rom[198][22] = 16'hFFEA;
        rom[198][23] = 16'hFFF4;
        rom[198][24] = 16'hFFF3;
        rom[198][25] = 16'h000A;
        rom[198][26] = 16'hFFDC;
        rom[198][27] = 16'hFFF9;
        rom[198][28] = 16'hFFDD;
        rom[198][29] = 16'h0016;
        rom[198][30] = 16'h0010;
        rom[198][31] = 16'h0044;
        rom[198][32] = 16'hFFE5;
        rom[198][33] = 16'h0004;
        rom[198][34] = 16'h003A;
        rom[198][35] = 16'h001A;
        rom[198][36] = 16'hFFF9;
        rom[198][37] = 16'hFFE5;
        rom[198][38] = 16'h005A;
        rom[198][39] = 16'h0028;
        rom[198][40] = 16'hFFF9;
        rom[198][41] = 16'h002E;
        rom[198][42] = 16'hFFF1;
        rom[198][43] = 16'h0006;
        rom[198][44] = 16'h0035;
        rom[198][45] = 16'hFFF5;
        rom[198][46] = 16'h000A;
        rom[198][47] = 16'hFFFE;
        rom[198][48] = 16'hFFD8;
        rom[198][49] = 16'hFFC5;
        rom[198][50] = 16'h001D;
        rom[198][51] = 16'hFFFD;
        rom[198][52] = 16'h0002;
        rom[198][53] = 16'hFFCB;
        rom[198][54] = 16'h001E;
        rom[198][55] = 16'h0028;
        rom[198][56] = 16'hFFE6;
        rom[198][57] = 16'h000D;
        rom[198][58] = 16'h000C;
        rom[198][59] = 16'hFFEE;
        rom[198][60] = 16'hFFF1;
        rom[198][61] = 16'h0002;
        rom[198][62] = 16'h0007;
        rom[198][63] = 16'h001F;
        rom[198][64] = 16'hFFFC;
        rom[198][65] = 16'hFFFD;
        rom[198][66] = 16'hFFE0;
        rom[198][67] = 16'hFFEA;
        rom[198][68] = 16'hFFDC;
        rom[198][69] = 16'hFFF3;
        rom[198][70] = 16'h000E;
        rom[198][71] = 16'hFFE0;
        rom[198][72] = 16'h0004;
        rom[198][73] = 16'h001F;
        rom[198][74] = 16'h001B;
        rom[198][75] = 16'h0026;
        rom[198][76] = 16'h001A;
        rom[198][77] = 16'hFFF1;
        rom[198][78] = 16'hFFEE;
        rom[198][79] = 16'h0016;
        rom[198][80] = 16'hFFD4;
        rom[198][81] = 16'h0002;
        rom[198][82] = 16'hFFD8;
        rom[198][83] = 16'h0016;
        rom[198][84] = 16'h0016;
        rom[198][85] = 16'hFFEA;
        rom[198][86] = 16'hFFE0;
        rom[198][87] = 16'hFFFA;
        rom[198][88] = 16'hFFEA;
        rom[198][89] = 16'hFFFD;
        rom[198][90] = 16'hFFE8;
        rom[198][91] = 16'hFFD4;
        rom[198][92] = 16'h0007;
        rom[198][93] = 16'h0016;
        rom[198][94] = 16'hFFE9;
        rom[198][95] = 16'hFFAD;
        rom[198][96] = 16'hFFE9;
        rom[198][97] = 16'h000B;
        rom[198][98] = 16'h0000;
        rom[198][99] = 16'hFFC8;
        rom[198][100] = 16'hFFEE;
        rom[198][101] = 16'h0014;
        rom[198][102] = 16'hFFF0;
        rom[198][103] = 16'hFFEF;
        rom[198][104] = 16'hFFFE;
        rom[198][105] = 16'hFFED;
        rom[198][106] = 16'hFFF9;
        rom[198][107] = 16'hFFF1;
        rom[198][108] = 16'hFFBD;
        rom[198][109] = 16'hFFF3;
        rom[198][110] = 16'hFFD6;
        rom[198][111] = 16'hFFCF;
        rom[198][112] = 16'hFFEA;
        rom[198][113] = 16'h0002;
        rom[198][114] = 16'hFFEE;
        rom[198][115] = 16'h0012;
        rom[198][116] = 16'h0020;
        rom[198][117] = 16'hFFF1;
        rom[198][118] = 16'hFFCD;
        rom[198][119] = 16'h0023;
        rom[198][120] = 16'hFFD8;
        rom[198][121] = 16'hFFE8;
        rom[198][122] = 16'h0028;
        rom[198][123] = 16'h0020;
        rom[198][124] = 16'h0004;
        rom[198][125] = 16'h001A;
        rom[198][126] = 16'hFFC8;
        rom[198][127] = 16'h0008;
        rom[199][0] = 16'hFFC8;
        rom[199][1] = 16'h000C;
        rom[199][2] = 16'h0015;
        rom[199][3] = 16'h000D;
        rom[199][4] = 16'h0002;
        rom[199][5] = 16'h0012;
        rom[199][6] = 16'hFFCE;
        rom[199][7] = 16'hFFF3;
        rom[199][8] = 16'h0001;
        rom[199][9] = 16'hFFB2;
        rom[199][10] = 16'hFFE5;
        rom[199][11] = 16'hFFB0;
        rom[199][12] = 16'hFFEA;
        rom[199][13] = 16'h0009;
        rom[199][14] = 16'hFFE7;
        rom[199][15] = 16'h0007;
        rom[199][16] = 16'h000C;
        rom[199][17] = 16'h000C;
        rom[199][18] = 16'hFFCD;
        rom[199][19] = 16'hFFEA;
        rom[199][20] = 16'hFFD0;
        rom[199][21] = 16'h0033;
        rom[199][22] = 16'hFFCB;
        rom[199][23] = 16'hFFD0;
        rom[199][24] = 16'hFFC3;
        rom[199][25] = 16'hFFEE;
        rom[199][26] = 16'hFFF1;
        rom[199][27] = 16'h003C;
        rom[199][28] = 16'h0005;
        rom[199][29] = 16'h0014;
        rom[199][30] = 16'h001B;
        rom[199][31] = 16'hFFDC;
        rom[199][32] = 16'hFFFF;
        rom[199][33] = 16'hFFEA;
        rom[199][34] = 16'h0002;
        rom[199][35] = 16'h0019;
        rom[199][36] = 16'hFFDB;
        rom[199][37] = 16'hFFEF;
        rom[199][38] = 16'hFFCE;
        rom[199][39] = 16'h0006;
        rom[199][40] = 16'hFFCF;
        rom[199][41] = 16'hFFC9;
        rom[199][42] = 16'hFFF4;
        rom[199][43] = 16'h001A;
        rom[199][44] = 16'h0016;
        rom[199][45] = 16'h0002;
        rom[199][46] = 16'hFFD3;
        rom[199][47] = 16'hFFF9;
        rom[199][48] = 16'hFFF7;
        rom[199][49] = 16'h0026;
        rom[199][50] = 16'hFFDC;
        rom[199][51] = 16'h0005;
        rom[199][52] = 16'h0025;
        rom[199][53] = 16'h0006;
        rom[199][54] = 16'h0021;
        rom[199][55] = 16'h000E;
        rom[199][56] = 16'h0009;
        rom[199][57] = 16'h0002;
        rom[199][58] = 16'h001C;
        rom[199][59] = 16'hFFE4;
        rom[199][60] = 16'hFFF5;
        rom[199][61] = 16'h0006;
        rom[199][62] = 16'hFFE6;
        rom[199][63] = 16'hFFF7;
        rom[199][64] = 16'hFFFF;
        rom[199][65] = 16'hFFD2;
        rom[199][66] = 16'h0005;
        rom[199][67] = 16'h0013;
        rom[199][68] = 16'hFFF1;
        rom[199][69] = 16'h0001;
        rom[199][70] = 16'hFFED;
        rom[199][71] = 16'h0011;
        rom[199][72] = 16'hFFDC;
        rom[199][73] = 16'hFFF9;
        rom[199][74] = 16'hFFCD;
        rom[199][75] = 16'hFFC8;
        rom[199][76] = 16'hFFD2;
        rom[199][77] = 16'h0037;
        rom[199][78] = 16'hFFE1;
        rom[199][79] = 16'h001E;
        rom[199][80] = 16'h001C;
        rom[199][81] = 16'hFFFA;
        rom[199][82] = 16'h0007;
        rom[199][83] = 16'h0000;
        rom[199][84] = 16'h000B;
        rom[199][85] = 16'hFFFB;
        rom[199][86] = 16'hFFDB;
        rom[199][87] = 16'hFFF4;
        rom[199][88] = 16'hFFBC;
        rom[199][89] = 16'h002A;
        rom[199][90] = 16'hFFF1;
        rom[199][91] = 16'hFFFF;
        rom[199][92] = 16'hFFC4;
        rom[199][93] = 16'h000E;
        rom[199][94] = 16'hFFE8;
        rom[199][95] = 16'hFF9D;
        rom[199][96] = 16'h0017;
        rom[199][97] = 16'hFFD3;
        rom[199][98] = 16'h000C;
        rom[199][99] = 16'h000E;
        rom[199][100] = 16'hFFE9;
        rom[199][101] = 16'h0005;
        rom[199][102] = 16'hFFCC;
        rom[199][103] = 16'h0019;
        rom[199][104] = 16'h0032;
        rom[199][105] = 16'h000C;
        rom[199][106] = 16'hFFFD;
        rom[199][107] = 16'h000E;
        rom[199][108] = 16'hFFF7;
        rom[199][109] = 16'hFFEF;
        rom[199][110] = 16'h0002;
        rom[199][111] = 16'hFFEF;
        rom[199][112] = 16'hFFE1;
        rom[199][113] = 16'hFFD9;
        rom[199][114] = 16'h004D;
        rom[199][115] = 16'hFFF3;
        rom[199][116] = 16'hFFD8;
        rom[199][117] = 16'hFFE1;
        rom[199][118] = 16'hFFBF;
        rom[199][119] = 16'hFFDB;
        rom[199][120] = 16'hFFD1;
        rom[199][121] = 16'hFFEA;
        rom[199][122] = 16'hFFF0;
        rom[199][123] = 16'hFFE1;
        rom[199][124] = 16'h0019;
        rom[199][125] = 16'hFFF0;
        rom[199][126] = 16'h0022;
        rom[199][127] = 16'h000F;
        rom[200][0] = 16'hFFD7;
        rom[200][1] = 16'h000C;
        rom[200][2] = 16'h002E;
        rom[200][3] = 16'hFFDB;
        rom[200][4] = 16'hFFEF;
        rom[200][5] = 16'h000E;
        rom[200][6] = 16'hFFF3;
        rom[200][7] = 16'h001B;
        rom[200][8] = 16'hFFF4;
        rom[200][9] = 16'h0025;
        rom[200][10] = 16'hFFF4;
        rom[200][11] = 16'hFFDA;
        rom[200][12] = 16'h0001;
        rom[200][13] = 16'h0002;
        rom[200][14] = 16'h001B;
        rom[200][15] = 16'h0013;
        rom[200][16] = 16'hFFC9;
        rom[200][17] = 16'hFFEA;
        rom[200][18] = 16'h0012;
        rom[200][19] = 16'h0013;
        rom[200][20] = 16'hFFD5;
        rom[200][21] = 16'h0019;
        rom[200][22] = 16'h000C;
        rom[200][23] = 16'h000F;
        rom[200][24] = 16'h0017;
        rom[200][25] = 16'h000C;
        rom[200][26] = 16'h0008;
        rom[200][27] = 16'hFFBC;
        rom[200][28] = 16'hFFD8;
        rom[200][29] = 16'hFFF7;
        rom[200][30] = 16'hFFF4;
        rom[200][31] = 16'h001C;
        rom[200][32] = 16'h001E;
        rom[200][33] = 16'h0012;
        rom[200][34] = 16'hFFFD;
        rom[200][35] = 16'h001F;
        rom[200][36] = 16'h000C;
        rom[200][37] = 16'hFFEF;
        rom[200][38] = 16'hFFF1;
        rom[200][39] = 16'hFFFA;
        rom[200][40] = 16'hFFF0;
        rom[200][41] = 16'hFFF8;
        rom[200][42] = 16'hFFFD;
        rom[200][43] = 16'hFFCC;
        rom[200][44] = 16'h000C;
        rom[200][45] = 16'h002E;
        rom[200][46] = 16'h0002;
        rom[200][47] = 16'h0028;
        rom[200][48] = 16'h0011;
        rom[200][49] = 16'h0011;
        rom[200][50] = 16'h0011;
        rom[200][51] = 16'hFFC8;
        rom[200][52] = 16'hFFC7;
        rom[200][53] = 16'hFFFA;
        rom[200][54] = 16'h000C;
        rom[200][55] = 16'hFFF4;
        rom[200][56] = 16'hFFFD;
        rom[200][57] = 16'hFFCE;
        rom[200][58] = 16'h0007;
        rom[200][59] = 16'hFFE1;
        rom[200][60] = 16'hFFFB;
        rom[200][61] = 16'h0011;
        rom[200][62] = 16'h0025;
        rom[200][63] = 16'h000C;
        rom[200][64] = 16'hFFE6;
        rom[200][65] = 16'hFFFF;
        rom[200][66] = 16'h0023;
        rom[200][67] = 16'h0002;
        rom[200][68] = 16'hFFFE;
        rom[200][69] = 16'h000C;
        rom[200][70] = 16'h003C;
        rom[200][71] = 16'hFFD4;
        rom[200][72] = 16'h0000;
        rom[200][73] = 16'h000A;
        rom[200][74] = 16'hFFF9;
        rom[200][75] = 16'h0016;
        rom[200][76] = 16'hFFEB;
        rom[200][77] = 16'hFFD0;
        rom[200][78] = 16'hFFEF;
        rom[200][79] = 16'h0002;
        rom[200][80] = 16'h001E;
        rom[200][81] = 16'h001A;
        rom[200][82] = 16'h0010;
        rom[200][83] = 16'hFFFB;
        rom[200][84] = 16'hFFF1;
        rom[200][85] = 16'hFFF3;
        rom[200][86] = 16'h001B;
        rom[200][87] = 16'hFF9C;
        rom[200][88] = 16'hFFD1;
        rom[200][89] = 16'h0009;
        rom[200][90] = 16'h0009;
        rom[200][91] = 16'hFFB0;
        rom[200][92] = 16'h0008;
        rom[200][93] = 16'h0010;
        rom[200][94] = 16'hFFD2;
        rom[200][95] = 16'hFFCB;
        rom[200][96] = 16'hFFB2;
        rom[200][97] = 16'hFFBA;
        rom[200][98] = 16'hFFB5;
        rom[200][99] = 16'h000C;
        rom[200][100] = 16'hFFA6;
        rom[200][101] = 16'h0002;
        rom[200][102] = 16'hFFF8;
        rom[200][103] = 16'hFFB5;
        rom[200][104] = 16'hFFD2;
        rom[200][105] = 16'hFFC8;
        rom[200][106] = 16'hFFEF;
        rom[200][107] = 16'h0027;
        rom[200][108] = 16'hFFCC;
        rom[200][109] = 16'hFFF9;
        rom[200][110] = 16'hFFFB;
        rom[200][111] = 16'hFFE8;
        rom[200][112] = 16'hFFE8;
        rom[200][113] = 16'hFFCC;
        rom[200][114] = 16'hFFFC;
        rom[200][115] = 16'h0038;
        rom[200][116] = 16'hFFEF;
        rom[200][117] = 16'h0026;
        rom[200][118] = 16'h0012;
        rom[200][119] = 16'h0025;
        rom[200][120] = 16'hFFE1;
        rom[200][121] = 16'h0018;
        rom[200][122] = 16'hFFF8;
        rom[200][123] = 16'hFFF9;
        rom[200][124] = 16'h0010;
        rom[200][125] = 16'hFFBA;
        rom[200][126] = 16'hFFB8;
        rom[200][127] = 16'hFFF1;
        rom[201][0] = 16'h000E;
        rom[201][1] = 16'h0016;
        rom[201][2] = 16'h0027;
        rom[201][3] = 16'h0027;
        rom[201][4] = 16'hFFDA;
        rom[201][5] = 16'hFFF9;
        rom[201][6] = 16'h0007;
        rom[201][7] = 16'hFFFF;
        rom[201][8] = 16'h0011;
        rom[201][9] = 16'h001D;
        rom[201][10] = 16'h0002;
        rom[201][11] = 16'hFFFA;
        rom[201][12] = 16'h0013;
        rom[201][13] = 16'hFFEA;
        rom[201][14] = 16'h003D;
        rom[201][15] = 16'hFFEE;
        rom[201][16] = 16'hFFF4;
        rom[201][17] = 16'h000A;
        rom[201][18] = 16'hFFFA;
        rom[201][19] = 16'h0011;
        rom[201][20] = 16'hFFDB;
        rom[201][21] = 16'h0016;
        rom[201][22] = 16'h000F;
        rom[201][23] = 16'hFFE9;
        rom[201][24] = 16'h0012;
        rom[201][25] = 16'hFFB6;
        rom[201][26] = 16'h0027;
        rom[201][27] = 16'hFFEA;
        rom[201][28] = 16'h0007;
        rom[201][29] = 16'h0010;
        rom[201][30] = 16'hFFFC;
        rom[201][31] = 16'hFFD7;
        rom[201][32] = 16'h001B;
        rom[201][33] = 16'h001A;
        rom[201][34] = 16'hFFEA;
        rom[201][35] = 16'h001A;
        rom[201][36] = 16'hFFEF;
        rom[201][37] = 16'h0011;
        rom[201][38] = 16'h000F;
        rom[201][39] = 16'h0018;
        rom[201][40] = 16'hFFF3;
        rom[201][41] = 16'h0004;
        rom[201][42] = 16'h0017;
        rom[201][43] = 16'hFFD3;
        rom[201][44] = 16'hFFD3;
        rom[201][45] = 16'h0025;
        rom[201][46] = 16'hFFEA;
        rom[201][47] = 16'hFFF0;
        rom[201][48] = 16'h0023;
        rom[201][49] = 16'h001B;
        rom[201][50] = 16'h000E;
        rom[201][51] = 16'hFFE8;
        rom[201][52] = 16'hFFEB;
        rom[201][53] = 16'h0017;
        rom[201][54] = 16'hFFE0;
        rom[201][55] = 16'hFFAA;
        rom[201][56] = 16'h0002;
        rom[201][57] = 16'h0006;
        rom[201][58] = 16'hFFF9;
        rom[201][59] = 16'hFFE2;
        rom[201][60] = 16'hFFB5;
        rom[201][61] = 16'hFFEF;
        rom[201][62] = 16'hFFE7;
        rom[201][63] = 16'hFFC5;
        rom[201][64] = 16'h0016;
        rom[201][65] = 16'h000B;
        rom[201][66] = 16'h0016;
        rom[201][67] = 16'h000C;
        rom[201][68] = 16'hFFE4;
        rom[201][69] = 16'hFFEA;
        rom[201][70] = 16'h0029;
        rom[201][71] = 16'h0033;
        rom[201][72] = 16'hFFEA;
        rom[201][73] = 16'hFFE9;
        rom[201][74] = 16'hFFDD;
        rom[201][75] = 16'h0024;
        rom[201][76] = 16'h000E;
        rom[201][77] = 16'hFFDC;
        rom[201][78] = 16'hFFF3;
        rom[201][79] = 16'h0017;
        rom[201][80] = 16'h000D;
        rom[201][81] = 16'hFFEF;
        rom[201][82] = 16'h000A;
        rom[201][83] = 16'h001B;
        rom[201][84] = 16'h001F;
        rom[201][85] = 16'hFFE5;
        rom[201][86] = 16'h0009;
        rom[201][87] = 16'hFFC5;
        rom[201][88] = 16'hFFC0;
        rom[201][89] = 16'hFFF4;
        rom[201][90] = 16'hFFEF;
        rom[201][91] = 16'h0024;
        rom[201][92] = 16'h000A;
        rom[201][93] = 16'h000A;
        rom[201][94] = 16'hFFCB;
        rom[201][95] = 16'hFFD7;
        rom[201][96] = 16'hFFF0;
        rom[201][97] = 16'h0004;
        rom[201][98] = 16'hFFEC;
        rom[201][99] = 16'hFFC3;
        rom[201][100] = 16'hFFF5;
        rom[201][101] = 16'hFFFC;
        rom[201][102] = 16'hFFFE;
        rom[201][103] = 16'h0008;
        rom[201][104] = 16'hFFEE;
        rom[201][105] = 16'h0021;
        rom[201][106] = 16'hFFFD;
        rom[201][107] = 16'h0006;
        rom[201][108] = 16'hFFFB;
        rom[201][109] = 16'hFFF8;
        rom[201][110] = 16'h0027;
        rom[201][111] = 16'hFFD7;
        rom[201][112] = 16'h0001;
        rom[201][113] = 16'hFFD5;
        rom[201][114] = 16'h0018;
        rom[201][115] = 16'hFFE7;
        rom[201][116] = 16'hFFEB;
        rom[201][117] = 16'h001F;
        rom[201][118] = 16'hFFEF;
        rom[201][119] = 16'h0021;
        rom[201][120] = 16'hFFD7;
        rom[201][121] = 16'hFFFB;
        rom[201][122] = 16'hFFF0;
        rom[201][123] = 16'hFFDB;
        rom[201][124] = 16'hFFE8;
        rom[201][125] = 16'hFFE7;
        rom[201][126] = 16'hFFF8;
        rom[201][127] = 16'hFFFE;
        rom[202][0] = 16'h0030;
        rom[202][1] = 16'h0024;
        rom[202][2] = 16'hFFDA;
        rom[202][3] = 16'hFFCC;
        rom[202][4] = 16'h0025;
        rom[202][5] = 16'h000A;
        rom[202][6] = 16'h0010;
        rom[202][7] = 16'hFFF3;
        rom[202][8] = 16'h003F;
        rom[202][9] = 16'hFFBA;
        rom[202][10] = 16'hFFBF;
        rom[202][11] = 16'h0002;
        rom[202][12] = 16'hFFE2;
        rom[202][13] = 16'h0011;
        rom[202][14] = 16'hFFE4;
        rom[202][15] = 16'hFFB1;
        rom[202][16] = 16'hFFFA;
        rom[202][17] = 16'h000F;
        rom[202][18] = 16'h002C;
        rom[202][19] = 16'h0024;
        rom[202][20] = 16'h0018;
        rom[202][21] = 16'hFFD7;
        rom[202][22] = 16'h0019;
        rom[202][23] = 16'h0016;
        rom[202][24] = 16'hFFE4;
        rom[202][25] = 16'h0007;
        rom[202][26] = 16'h0032;
        rom[202][27] = 16'hFFDE;
        rom[202][28] = 16'hFFE5;
        rom[202][29] = 16'h0006;
        rom[202][30] = 16'h0026;
        rom[202][31] = 16'h0007;
        rom[202][32] = 16'h0003;
        rom[202][33] = 16'hFFE4;
        rom[202][34] = 16'hFFF4;
        rom[202][35] = 16'hFFC7;
        rom[202][36] = 16'hFFF7;
        rom[202][37] = 16'h0024;
        rom[202][38] = 16'hFFD2;
        rom[202][39] = 16'hFFF9;
        rom[202][40] = 16'h0007;
        rom[202][41] = 16'h0009;
        rom[202][42] = 16'hFFDD;
        rom[202][43] = 16'hFFE8;
        rom[202][44] = 16'hFFEC;
        rom[202][45] = 16'hFFB8;
        rom[202][46] = 16'hFFE6;
        rom[202][47] = 16'h0006;
        rom[202][48] = 16'hFFEA;
        rom[202][49] = 16'h0028;
        rom[202][50] = 16'hFFD0;
        rom[202][51] = 16'h0021;
        rom[202][52] = 16'hFFFE;
        rom[202][53] = 16'hFFDF;
        rom[202][54] = 16'hFFBF;
        rom[202][55] = 16'hFFF3;
        rom[202][56] = 16'h000C;
        rom[202][57] = 16'h003B;
        rom[202][58] = 16'hFFCE;
        rom[202][59] = 16'h0006;
        rom[202][60] = 16'hFFBF;
        rom[202][61] = 16'hFFF9;
        rom[202][62] = 16'hFFFA;
        rom[202][63] = 16'h001A;
        rom[202][64] = 16'h000E;
        rom[202][65] = 16'h0000;
        rom[202][66] = 16'h0006;
        rom[202][67] = 16'h0025;
        rom[202][68] = 16'hFFEA;
        rom[202][69] = 16'hFFE5;
        rom[202][70] = 16'hFFD3;
        rom[202][71] = 16'h0024;
        rom[202][72] = 16'h002F;
        rom[202][73] = 16'h0016;
        rom[202][74] = 16'h0004;
        rom[202][75] = 16'hFFD8;
        rom[202][76] = 16'hFFE7;
        rom[202][77] = 16'hFFB8;
        rom[202][78] = 16'h0025;
        rom[202][79] = 16'h0002;
        rom[202][80] = 16'hFFEA;
        rom[202][81] = 16'h000C;
        rom[202][82] = 16'h0033;
        rom[202][83] = 16'hFFE7;
        rom[202][84] = 16'hFFE2;
        rom[202][85] = 16'hFFB7;
        rom[202][86] = 16'h0018;
        rom[202][87] = 16'h0040;
        rom[202][88] = 16'h000E;
        rom[202][89] = 16'hFFCF;
        rom[202][90] = 16'h0038;
        rom[202][91] = 16'h000A;
        rom[202][92] = 16'hFFFD;
        rom[202][93] = 16'hFFFB;
        rom[202][94] = 16'hFFFB;
        rom[202][95] = 16'h0015;
        rom[202][96] = 16'hFFF9;
        rom[202][97] = 16'h001F;
        rom[202][98] = 16'h0017;
        rom[202][99] = 16'hFFFE;
        rom[202][100] = 16'h000A;
        rom[202][101] = 16'h001D;
        rom[202][102] = 16'h0009;
        rom[202][103] = 16'h001C;
        rom[202][104] = 16'h0007;
        rom[202][105] = 16'h0029;
        rom[202][106] = 16'hFFEB;
        rom[202][107] = 16'hFF9C;
        rom[202][108] = 16'h001F;
        rom[202][109] = 16'hFFE6;
        rom[202][110] = 16'h0002;
        rom[202][111] = 16'hFFEF;
        rom[202][112] = 16'h000F;
        rom[202][113] = 16'h0006;
        rom[202][114] = 16'hFFF8;
        rom[202][115] = 16'hFFDD;
        rom[202][116] = 16'h0022;
        rom[202][117] = 16'hFFFC;
        rom[202][118] = 16'hFFEA;
        rom[202][119] = 16'hFFF7;
        rom[202][120] = 16'h0033;
        rom[202][121] = 16'hFFDE;
        rom[202][122] = 16'h001D;
        rom[202][123] = 16'hFFE7;
        rom[202][124] = 16'hFFDA;
        rom[202][125] = 16'h001A;
        rom[202][126] = 16'hFFC4;
        rom[202][127] = 16'hFFEF;
        rom[203][0] = 16'hFFDC;
        rom[203][1] = 16'hFFEA;
        rom[203][2] = 16'h0024;
        rom[203][3] = 16'hFFA4;
        rom[203][4] = 16'hFFE5;
        rom[203][5] = 16'hFFE7;
        rom[203][6] = 16'h000E;
        rom[203][7] = 16'hFFC6;
        rom[203][8] = 16'hFFD4;
        rom[203][9] = 16'hFFFB;
        rom[203][10] = 16'h0029;
        rom[203][11] = 16'h000C;
        rom[203][12] = 16'h0029;
        rom[203][13] = 16'hFFEF;
        rom[203][14] = 16'hFFE3;
        rom[203][15] = 16'h0013;
        rom[203][16] = 16'h0019;
        rom[203][17] = 16'hFFC9;
        rom[203][18] = 16'h0002;
        rom[203][19] = 16'h0001;
        rom[203][20] = 16'hFFB8;
        rom[203][21] = 16'hFFE7;
        rom[203][22] = 16'hFFDE;
        rom[203][23] = 16'hFFE3;
        rom[203][24] = 16'h000F;
        rom[203][25] = 16'h0011;
        rom[203][26] = 16'hFFFE;
        rom[203][27] = 16'hFFD6;
        rom[203][28] = 16'hFFE8;
        rom[203][29] = 16'h0025;
        rom[203][30] = 16'hFFD1;
        rom[203][31] = 16'hFFBE;
        rom[203][32] = 16'hFFEE;
        rom[203][33] = 16'h0009;
        rom[203][34] = 16'hFFE3;
        rom[203][35] = 16'hFFFD;
        rom[203][36] = 16'h0009;
        rom[203][37] = 16'h0001;
        rom[203][38] = 16'hFFE1;
        rom[203][39] = 16'h000E;
        rom[203][40] = 16'hFFF6;
        rom[203][41] = 16'hFFE9;
        rom[203][42] = 16'h0006;
        rom[203][43] = 16'h0001;
        rom[203][44] = 16'h0008;
        rom[203][45] = 16'hFFF6;
        rom[203][46] = 16'h0009;
        rom[203][47] = 16'hFFD4;
        rom[203][48] = 16'h0012;
        rom[203][49] = 16'h0024;
        rom[203][50] = 16'hFFFD;
        rom[203][51] = 16'hFFD8;
        rom[203][52] = 16'h0010;
        rom[203][53] = 16'h0009;
        rom[203][54] = 16'hFFCA;
        rom[203][55] = 16'h0000;
        rom[203][56] = 16'h001C;
        rom[203][57] = 16'hFFEB;
        rom[203][58] = 16'h0002;
        rom[203][59] = 16'h0005;
        rom[203][60] = 16'hFFE3;
        rom[203][61] = 16'h001A;
        rom[203][62] = 16'hFFCA;
        rom[203][63] = 16'hFFD3;
        rom[203][64] = 16'hFFDD;
        rom[203][65] = 16'hFFD0;
        rom[203][66] = 16'hFFF4;
        rom[203][67] = 16'h002F;
        rom[203][68] = 16'h000B;
        rom[203][69] = 16'h002E;
        rom[203][70] = 16'h0015;
        rom[203][71] = 16'h0009;
        rom[203][72] = 16'hFFDD;
        rom[203][73] = 16'h0030;
        rom[203][74] = 16'hFFB4;
        rom[203][75] = 16'h001D;
        rom[203][76] = 16'h0015;
        rom[203][77] = 16'h0018;
        rom[203][78] = 16'hFFD2;
        rom[203][79] = 16'h0007;
        rom[203][80] = 16'hFFCD;
        rom[203][81] = 16'hFFEA;
        rom[203][82] = 16'hFFEB;
        rom[203][83] = 16'h0020;
        rom[203][84] = 16'h0011;
        rom[203][85] = 16'h0006;
        rom[203][86] = 16'hFFF3;
        rom[203][87] = 16'hFFDC;
        rom[203][88] = 16'hFFB3;
        rom[203][89] = 16'hFFE1;
        rom[203][90] = 16'hFFE6;
        rom[203][91] = 16'hFFD6;
        rom[203][92] = 16'h000A;
        rom[203][93] = 16'hFFD0;
        rom[203][94] = 16'hFFF4;
        rom[203][95] = 16'hFFD2;
        rom[203][96] = 16'hFFB5;
        rom[203][97] = 16'hFFF2;
        rom[203][98] = 16'h0050;
        rom[203][99] = 16'h001A;
        rom[203][100] = 16'h0001;
        rom[203][101] = 16'hFFF8;
        rom[203][102] = 16'hFFDF;
        rom[203][103] = 16'hFFBC;
        rom[203][104] = 16'h0029;
        rom[203][105] = 16'hFFF2;
        rom[203][106] = 16'hFFF8;
        rom[203][107] = 16'h0033;
        rom[203][108] = 16'h0026;
        rom[203][109] = 16'hFFD2;
        rom[203][110] = 16'hFFE3;
        rom[203][111] = 16'h001D;
        rom[203][112] = 16'hFFFF;
        rom[203][113] = 16'hFFFF;
        rom[203][114] = 16'h0002;
        rom[203][115] = 16'hFFE7;
        rom[203][116] = 16'hFFCE;
        rom[203][117] = 16'hFFF8;
        rom[203][118] = 16'hFFCF;
        rom[203][119] = 16'hFFF2;
        rom[203][120] = 16'h0011;
        rom[203][121] = 16'hFFC8;
        rom[203][122] = 16'h003A;
        rom[203][123] = 16'hFFE9;
        rom[203][124] = 16'hFFEC;
        rom[203][125] = 16'hFFF1;
        rom[203][126] = 16'hFFF4;
        rom[203][127] = 16'h0032;
        rom[204][0] = 16'hFFFF;
        rom[204][1] = 16'hFFFA;
        rom[204][2] = 16'hFFF4;
        rom[204][3] = 16'h0028;
        rom[204][4] = 16'hFFD2;
        rom[204][5] = 16'hFFFB;
        rom[204][6] = 16'hFFF8;
        rom[204][7] = 16'hFFFF;
        rom[204][8] = 16'hFFC8;
        rom[204][9] = 16'h001F;
        rom[204][10] = 16'h0003;
        rom[204][11] = 16'hFFD2;
        rom[204][12] = 16'hFFD7;
        rom[204][13] = 16'hFFFE;
        rom[204][14] = 16'h0004;
        rom[204][15] = 16'h000C;
        rom[204][16] = 16'hFFE5;
        rom[204][17] = 16'hFFDE;
        rom[204][18] = 16'h000F;
        rom[204][19] = 16'h000C;
        rom[204][20] = 16'h0009;
        rom[204][21] = 16'h000F;
        rom[204][22] = 16'h0006;
        rom[204][23] = 16'h0007;
        rom[204][24] = 16'hFFF5;
        rom[204][25] = 16'h003D;
        rom[204][26] = 16'hFFFF;
        rom[204][27] = 16'h001E;
        rom[204][28] = 16'h0016;
        rom[204][29] = 16'h0001;
        rom[204][30] = 16'h0004;
        rom[204][31] = 16'h001B;
        rom[204][32] = 16'hFFDC;
        rom[204][33] = 16'h003C;
        rom[204][34] = 16'hFFD8;
        rom[204][35] = 16'h0010;
        rom[204][36] = 16'hFFD7;
        rom[204][37] = 16'hFFCC;
        rom[204][38] = 16'h0010;
        rom[204][39] = 16'hFFE6;
        rom[204][40] = 16'h001F;
        rom[204][41] = 16'h0011;
        rom[204][42] = 16'h0000;
        rom[204][43] = 16'hFFEC;
        rom[204][44] = 16'hFFEE;
        rom[204][45] = 16'h0011;
        rom[204][46] = 16'hFFC8;
        rom[204][47] = 16'h0004;
        rom[204][48] = 16'hFFE2;
        rom[204][49] = 16'hFFCC;
        rom[204][50] = 16'hFFE4;
        rom[204][51] = 16'h000E;
        rom[204][52] = 16'h0029;
        rom[204][53] = 16'hFFEC;
        rom[204][54] = 16'h0027;
        rom[204][55] = 16'h001C;
        rom[204][56] = 16'hFFE2;
        rom[204][57] = 16'hFFEC;
        rom[204][58] = 16'hFFF7;
        rom[204][59] = 16'hFFE1;
        rom[204][60] = 16'hFFFB;
        rom[204][61] = 16'hFFDA;
        rom[204][62] = 16'h000F;
        rom[204][63] = 16'h0012;
        rom[204][64] = 16'hFFDF;
        rom[204][65] = 16'h0013;
        rom[204][66] = 16'hFFEA;
        rom[204][67] = 16'h0007;
        rom[204][68] = 16'hFFEA;
        rom[204][69] = 16'hFFE5;
        rom[204][70] = 16'hFFFD;
        rom[204][71] = 16'h0014;
        rom[204][72] = 16'hFFD2;
        rom[204][73] = 16'h0007;
        rom[204][74] = 16'h0023;
        rom[204][75] = 16'h001F;
        rom[204][76] = 16'h000A;
        rom[204][77] = 16'hFFF6;
        rom[204][78] = 16'h002E;
        rom[204][79] = 16'h0007;
        rom[204][80] = 16'hFFFD;
        rom[204][81] = 16'h000D;
        rom[204][82] = 16'hFFE5;
        rom[204][83] = 16'hFFD2;
        rom[204][84] = 16'hFFF7;
        rom[204][85] = 16'hFFFB;
        rom[204][86] = 16'hFFFC;
        rom[204][87] = 16'h001B;
        rom[204][88] = 16'hFFDC;
        rom[204][89] = 16'h001F;
        rom[204][90] = 16'hFFDC;
        rom[204][91] = 16'h0001;
        rom[204][92] = 16'h002D;
        rom[204][93] = 16'h0009;
        rom[204][94] = 16'hFFD2;
        rom[204][95] = 16'h000C;
        rom[204][96] = 16'hFFFE;
        rom[204][97] = 16'hFFE4;
        rom[204][98] = 16'hFFC9;
        rom[204][99] = 16'hFFD9;
        rom[204][100] = 16'hFFF8;
        rom[204][101] = 16'h0025;
        rom[204][102] = 16'h0007;
        rom[204][103] = 16'h0020;
        rom[204][104] = 16'h0024;
        rom[204][105] = 16'h0027;
        rom[204][106] = 16'hFFCD;
        rom[204][107] = 16'hFFFE;
        rom[204][108] = 16'hFFE3;
        rom[204][109] = 16'h0016;
        rom[204][110] = 16'hFFCD;
        rom[204][111] = 16'h000C;
        rom[204][112] = 16'h0017;
        rom[204][113] = 16'hFFC3;
        rom[204][114] = 16'hFFDC;
        rom[204][115] = 16'hFFF9;
        rom[204][116] = 16'h0027;
        rom[204][117] = 16'hFFF5;
        rom[204][118] = 16'hFFEA;
        rom[204][119] = 16'h0027;
        rom[204][120] = 16'h0004;
        rom[204][121] = 16'hFFE8;
        rom[204][122] = 16'hFFE1;
        rom[204][123] = 16'h003C;
        rom[204][124] = 16'hFFF5;
        rom[204][125] = 16'h001A;
        rom[204][126] = 16'h0011;
        rom[204][127] = 16'h0005;
        rom[205][0] = 16'hFFFC;
        rom[205][1] = 16'h001B;
        rom[205][2] = 16'hFFE1;
        rom[205][3] = 16'h0013;
        rom[205][4] = 16'hFFD4;
        rom[205][5] = 16'hFFE2;
        rom[205][6] = 16'hFFFD;
        rom[205][7] = 16'h0011;
        rom[205][8] = 16'h0001;
        rom[205][9] = 16'hFFDA;
        rom[205][10] = 16'h000F;
        rom[205][11] = 16'h0006;
        rom[205][12] = 16'h0034;
        rom[205][13] = 16'hFFF8;
        rom[205][14] = 16'hFFDE;
        rom[205][15] = 16'hFFE1;
        rom[205][16] = 16'hFFF2;
        rom[205][17] = 16'h000D;
        rom[205][18] = 16'hFFCA;
        rom[205][19] = 16'h0022;
        rom[205][20] = 16'hFFD4;
        rom[205][21] = 16'h0012;
        rom[205][22] = 16'h000C;
        rom[205][23] = 16'h0021;
        rom[205][24] = 16'hFFEF;
        rom[205][25] = 16'h002B;
        rom[205][26] = 16'hFFE3;
        rom[205][27] = 16'h0031;
        rom[205][28] = 16'hFFE9;
        rom[205][29] = 16'hFFF4;
        rom[205][30] = 16'h0002;
        rom[205][31] = 16'h0011;
        rom[205][32] = 16'hFFE2;
        rom[205][33] = 16'h0001;
        rom[205][34] = 16'hFFF3;
        rom[205][35] = 16'h0024;
        rom[205][36] = 16'h0002;
        rom[205][37] = 16'hFFDD;
        rom[205][38] = 16'h0007;
        rom[205][39] = 16'h001B;
        rom[205][40] = 16'h0004;
        rom[205][41] = 16'hFFE0;
        rom[205][42] = 16'h0016;
        rom[205][43] = 16'hFFD4;
        rom[205][44] = 16'h001F;
        rom[205][45] = 16'h0032;
        rom[205][46] = 16'h000C;
        rom[205][47] = 16'h002A;
        rom[205][48] = 16'hFFE1;
        rom[205][49] = 16'hFFFA;
        rom[205][50] = 16'hFFF6;
        rom[205][51] = 16'h0002;
        rom[205][52] = 16'hFFFC;
        rom[205][53] = 16'h0008;
        rom[205][54] = 16'hFFEE;
        rom[205][55] = 16'hFFF9;
        rom[205][56] = 16'hFFD2;
        rom[205][57] = 16'h0004;
        rom[205][58] = 16'h0017;
        rom[205][59] = 16'h002B;
        rom[205][60] = 16'h0005;
        rom[205][61] = 16'h0038;
        rom[205][62] = 16'hFFF2;
        rom[205][63] = 16'hFFF6;
        rom[205][64] = 16'hFFE1;
        rom[205][65] = 16'hFFFC;
        rom[205][66] = 16'h000F;
        rom[205][67] = 16'hFFFD;
        rom[205][68] = 16'hFFDA;
        rom[205][69] = 16'h0036;
        rom[205][70] = 16'hFFF3;
        rom[205][71] = 16'hFFF7;
        rom[205][72] = 16'h0023;
        rom[205][73] = 16'hFFEF;
        rom[205][74] = 16'hFFF8;
        rom[205][75] = 16'h0011;
        rom[205][76] = 16'h0007;
        rom[205][77] = 16'h001F;
        rom[205][78] = 16'hFFF8;
        rom[205][79] = 16'h0014;
        rom[205][80] = 16'h001B;
        rom[205][81] = 16'h001A;
        rom[205][82] = 16'h0018;
        rom[205][83] = 16'h0023;
        rom[205][84] = 16'h0009;
        rom[205][85] = 16'hFFF9;
        rom[205][86] = 16'hFFE1;
        rom[205][87] = 16'h001B;
        rom[205][88] = 16'hFFFD;
        rom[205][89] = 16'hFFEB;
        rom[205][90] = 16'hFFFA;
        rom[205][91] = 16'h0010;
        rom[205][92] = 16'hFFFD;
        rom[205][93] = 16'h0019;
        rom[205][94] = 16'hFFD0;
        rom[205][95] = 16'hFFA6;
        rom[205][96] = 16'hFFE5;
        rom[205][97] = 16'hFFE5;
        rom[205][98] = 16'h0044;
        rom[205][99] = 16'h0022;
        rom[205][100] = 16'h0007;
        rom[205][101] = 16'h0006;
        rom[205][102] = 16'hFFE4;
        rom[205][103] = 16'h0014;
        rom[205][104] = 16'hFFF9;
        rom[205][105] = 16'hFFD2;
        rom[205][106] = 16'hFFDA;
        rom[205][107] = 16'h0029;
        rom[205][108] = 16'hFFBB;
        rom[205][109] = 16'hFFCD;
        rom[205][110] = 16'hFFDC;
        rom[205][111] = 16'h0028;
        rom[205][112] = 16'hFFE0;
        rom[205][113] = 16'hFFED;
        rom[205][114] = 16'h0011;
        rom[205][115] = 16'h000E;
        rom[205][116] = 16'h0023;
        rom[205][117] = 16'hFFE5;
        rom[205][118] = 16'hFFE6;
        rom[205][119] = 16'h001A;
        rom[205][120] = 16'h0006;
        rom[205][121] = 16'h000F;
        rom[205][122] = 16'h0029;
        rom[205][123] = 16'h0002;
        rom[205][124] = 16'hFFEE;
        rom[205][125] = 16'h0001;
        rom[205][126] = 16'hFFF4;
        rom[205][127] = 16'h0017;
        rom[206][0] = 16'h0020;
        rom[206][1] = 16'hFFAC;
        rom[206][2] = 16'hFFED;
        rom[206][3] = 16'h0013;
        rom[206][4] = 16'hFFE4;
        rom[206][5] = 16'hFFCC;
        rom[206][6] = 16'hFFDF;
        rom[206][7] = 16'hFFC8;
        rom[206][8] = 16'h0013;
        rom[206][9] = 16'h0015;
        rom[206][10] = 16'hFFE5;
        rom[206][11] = 16'h0006;
        rom[206][12] = 16'hFFE9;
        rom[206][13] = 16'h002C;
        rom[206][14] = 16'h001B;
        rom[206][15] = 16'h0011;
        rom[206][16] = 16'hFFCA;
        rom[206][17] = 16'hFFE5;
        rom[206][18] = 16'hFFFB;
        rom[206][19] = 16'h0012;
        rom[206][20] = 16'h000D;
        rom[206][21] = 16'hFFC3;
        rom[206][22] = 16'h001C;
        rom[206][23] = 16'hFFED;
        rom[206][24] = 16'h0006;
        rom[206][25] = 16'h0014;
        rom[206][26] = 16'hFFE1;
        rom[206][27] = 16'h000A;
        rom[206][28] = 16'hFFED;
        rom[206][29] = 16'h001C;
        rom[206][30] = 16'hFFD9;
        rom[206][31] = 16'h000C;
        rom[206][32] = 16'hFFEB;
        rom[206][33] = 16'hFFE6;
        rom[206][34] = 16'hFFD2;
        rom[206][35] = 16'hFFCD;
        rom[206][36] = 16'hFFBF;
        rom[206][37] = 16'hFFDA;
        rom[206][38] = 16'hFFED;
        rom[206][39] = 16'hFFE4;
        rom[206][40] = 16'hFFF8;
        rom[206][41] = 16'h000B;
        rom[206][42] = 16'hFFF6;
        rom[206][43] = 16'hFFEA;
        rom[206][44] = 16'hFFFB;
        rom[206][45] = 16'hFFD0;
        rom[206][46] = 16'hFFCD;
        rom[206][47] = 16'hFFFE;
        rom[206][48] = 16'hFFD4;
        rom[206][49] = 16'hFFC3;
        rom[206][50] = 16'hFFF9;
        rom[206][51] = 16'hFFED;
        rom[206][52] = 16'hFFF5;
        rom[206][53] = 16'hFFED;
        rom[206][54] = 16'hFFDF;
        rom[206][55] = 16'h0000;
        rom[206][56] = 16'hFFD8;
        rom[206][57] = 16'h000C;
        rom[206][58] = 16'hFFF6;
        rom[206][59] = 16'hFFE1;
        rom[206][60] = 16'h0002;
        rom[206][61] = 16'h0013;
        rom[206][62] = 16'hFFE9;
        rom[206][63] = 16'hFFE9;
        rom[206][64] = 16'hFFFF;
        rom[206][65] = 16'hFFF0;
        rom[206][66] = 16'h000C;
        rom[206][67] = 16'hFFF1;
        rom[206][68] = 16'hFFD7;
        rom[206][69] = 16'hFFE5;
        rom[206][70] = 16'hFFB9;
        rom[206][71] = 16'hFFF4;
        rom[206][72] = 16'hFFFD;
        rom[206][73] = 16'h0007;
        rom[206][74] = 16'hFFFE;
        rom[206][75] = 16'hFFEF;
        rom[206][76] = 16'hFFE2;
        rom[206][77] = 16'hFFE1;
        rom[206][78] = 16'h000D;
        rom[206][79] = 16'hFFD0;
        rom[206][80] = 16'h0009;
        rom[206][81] = 16'hFFD6;
        rom[206][82] = 16'hFFF0;
        rom[206][83] = 16'h001C;
        rom[206][84] = 16'hFFDB;
        rom[206][85] = 16'hFFFE;
        rom[206][86] = 16'hFFF3;
        rom[206][87] = 16'hFFD4;
        rom[206][88] = 16'hFFE9;
        rom[206][89] = 16'hFFEF;
        rom[206][90] = 16'h0007;
        rom[206][91] = 16'h0008;
        rom[206][92] = 16'h0026;
        rom[206][93] = 16'hFFC8;
        rom[206][94] = 16'h0016;
        rom[206][95] = 16'hFFF9;
        rom[206][96] = 16'hFFC3;
        rom[206][97] = 16'hFFC6;
        rom[206][98] = 16'hFFE7;
        rom[206][99] = 16'hFFE2;
        rom[206][100] = 16'hFFB8;
        rom[206][101] = 16'h001E;
        rom[206][102] = 16'hFFF8;
        rom[206][103] = 16'h0010;
        rom[206][104] = 16'hFFFE;
        rom[206][105] = 16'h002A;
        rom[206][106] = 16'h0012;
        rom[206][107] = 16'hFF9F;
        rom[206][108] = 16'hFFCF;
        rom[206][109] = 16'hFFDD;
        rom[206][110] = 16'hFFFE;
        rom[206][111] = 16'h0018;
        rom[206][112] = 16'h0011;
        rom[206][113] = 16'hFFF9;
        rom[206][114] = 16'hFFDA;
        rom[206][115] = 16'hFFD0;
        rom[206][116] = 16'hFFF4;
        rom[206][117] = 16'hFFFF;
        rom[206][118] = 16'hFFFF;
        rom[206][119] = 16'hFFD6;
        rom[206][120] = 16'h0025;
        rom[206][121] = 16'hFFFE;
        rom[206][122] = 16'hFFF3;
        rom[206][123] = 16'h001B;
        rom[206][124] = 16'hFFB5;
        rom[206][125] = 16'h000E;
        rom[206][126] = 16'hFFF2;
        rom[206][127] = 16'hFFCF;
        rom[207][0] = 16'hFFF4;
        rom[207][1] = 16'h0001;
        rom[207][2] = 16'hFFC5;
        rom[207][3] = 16'hFFD5;
        rom[207][4] = 16'h0004;
        rom[207][5] = 16'h001A;
        rom[207][6] = 16'hFFCD;
        rom[207][7] = 16'h0004;
        rom[207][8] = 16'h001B;
        rom[207][9] = 16'hFFDC;
        rom[207][10] = 16'h0024;
        rom[207][11] = 16'hFFD2;
        rom[207][12] = 16'hFFFD;
        rom[207][13] = 16'h0018;
        rom[207][14] = 16'h0016;
        rom[207][15] = 16'hFFED;
        rom[207][16] = 16'hFFEF;
        rom[207][17] = 16'h0010;
        rom[207][18] = 16'h001C;
        rom[207][19] = 16'hFFE6;
        rom[207][20] = 16'h0033;
        rom[207][21] = 16'h0022;
        rom[207][22] = 16'hFFF7;
        rom[207][23] = 16'h0024;
        rom[207][24] = 16'hFFF5;
        rom[207][25] = 16'h0021;
        rom[207][26] = 16'h0028;
        rom[207][27] = 16'h002B;
        rom[207][28] = 16'hFFCB;
        rom[207][29] = 16'hFFC2;
        rom[207][30] = 16'h0022;
        rom[207][31] = 16'h0024;
        rom[207][32] = 16'hFFD4;
        rom[207][33] = 16'h003F;
        rom[207][34] = 16'hFFC4;
        rom[207][35] = 16'hFFF9;
        rom[207][36] = 16'hFFE8;
        rom[207][37] = 16'hFFDB;
        rom[207][38] = 16'h000F;
        rom[207][39] = 16'hFFF4;
        rom[207][40] = 16'h000C;
        rom[207][41] = 16'h0015;
        rom[207][42] = 16'hFFFF;
        rom[207][43] = 16'hFFEC;
        rom[207][44] = 16'h000B;
        rom[207][45] = 16'hFFFE;
        rom[207][46] = 16'hFFF1;
        rom[207][47] = 16'hFFF4;
        rom[207][48] = 16'h0002;
        rom[207][49] = 16'h000B;
        rom[207][50] = 16'hFFAA;
        rom[207][51] = 16'h0029;
        rom[207][52] = 16'hFFAE;
        rom[207][53] = 16'h0035;
        rom[207][54] = 16'hFFDA;
        rom[207][55] = 16'hFFFE;
        rom[207][56] = 16'h000C;
        rom[207][57] = 16'h0003;
        rom[207][58] = 16'h0003;
        rom[207][59] = 16'h0011;
        rom[207][60] = 16'hFFFA;
        rom[207][61] = 16'hFFC4;
        rom[207][62] = 16'hFFEA;
        rom[207][63] = 16'h0002;
        rom[207][64] = 16'hFFF0;
        rom[207][65] = 16'h002B;
        rom[207][66] = 16'h0016;
        rom[207][67] = 16'h002A;
        rom[207][68] = 16'h0024;
        rom[207][69] = 16'h0012;
        rom[207][70] = 16'h0011;
        rom[207][71] = 16'hFFFE;
        rom[207][72] = 16'hFFFC;
        rom[207][73] = 16'h0027;
        rom[207][74] = 16'h000E;
        rom[207][75] = 16'h0014;
        rom[207][76] = 16'hFFF0;
        rom[207][77] = 16'hFFF1;
        rom[207][78] = 16'hFFE9;
        rom[207][79] = 16'hFFF4;
        rom[207][80] = 16'h0008;
        rom[207][81] = 16'hFFDD;
        rom[207][82] = 16'h0007;
        rom[207][83] = 16'h0016;
        rom[207][84] = 16'hFFFB;
        rom[207][85] = 16'hFFED;
        rom[207][86] = 16'hFFF6;
        rom[207][87] = 16'h000E;
        rom[207][88] = 16'h003D;
        rom[207][89] = 16'hFFFF;
        rom[207][90] = 16'h0024;
        rom[207][91] = 16'hFFFB;
        rom[207][92] = 16'h0019;
        rom[207][93] = 16'hFFEC;
        rom[207][94] = 16'h0002;
        rom[207][95] = 16'h000E;
        rom[207][96] = 16'h0000;
        rom[207][97] = 16'h0016;
        rom[207][98] = 16'h000A;
        rom[207][99] = 16'hFFE5;
        rom[207][100] = 16'hFFF9;
        rom[207][101] = 16'hFFD1;
        rom[207][102] = 16'hFFD9;
        rom[207][103] = 16'h0019;
        rom[207][104] = 16'h0018;
        rom[207][105] = 16'hFFD2;
        rom[207][106] = 16'hFFFC;
        rom[207][107] = 16'hFFE1;
        rom[207][108] = 16'hFFF1;
        rom[207][109] = 16'hFFF7;
        rom[207][110] = 16'hFFF8;
        rom[207][111] = 16'hFFEB;
        rom[207][112] = 16'h0024;
        rom[207][113] = 16'hFFFC;
        rom[207][114] = 16'h000B;
        rom[207][115] = 16'h0018;
        rom[207][116] = 16'hFFF6;
        rom[207][117] = 16'hFFEA;
        rom[207][118] = 16'hFFEA;
        rom[207][119] = 16'h0004;
        rom[207][120] = 16'hFFE7;
        rom[207][121] = 16'hFFD6;
        rom[207][122] = 16'hFFB2;
        rom[207][123] = 16'hFFE4;
        rom[207][124] = 16'hFFED;
        rom[207][125] = 16'h0009;
        rom[207][126] = 16'hFFE4;
        rom[207][127] = 16'hFFE8;
        rom[208][0] = 16'h0010;
        rom[208][1] = 16'hFFFD;
        rom[208][2] = 16'h0010;
        rom[208][3] = 16'hFFD9;
        rom[208][4] = 16'hFFF0;
        rom[208][5] = 16'h001B;
        rom[208][6] = 16'h0029;
        rom[208][7] = 16'hFFFA;
        rom[208][8] = 16'h001F;
        rom[208][9] = 16'h0017;
        rom[208][10] = 16'hFFCE;
        rom[208][11] = 16'hFFC1;
        rom[208][12] = 16'hFFDE;
        rom[208][13] = 16'h002E;
        rom[208][14] = 16'h000C;
        rom[208][15] = 16'h0016;
        rom[208][16] = 16'hFFEE;
        rom[208][17] = 16'hFFFF;
        rom[208][18] = 16'h0013;
        rom[208][19] = 16'h0024;
        rom[208][20] = 16'hFFEF;
        rom[208][21] = 16'h0001;
        rom[208][22] = 16'h0036;
        rom[208][23] = 16'hFFD2;
        rom[208][24] = 16'hFFF5;
        rom[208][25] = 16'hFFEF;
        rom[208][26] = 16'h000D;
        rom[208][27] = 16'h0014;
        rom[208][28] = 16'h0002;
        rom[208][29] = 16'h0024;
        rom[208][30] = 16'hFFBF;
        rom[208][31] = 16'h0029;
        rom[208][32] = 16'h0018;
        rom[208][33] = 16'h0007;
        rom[208][34] = 16'h0005;
        rom[208][35] = 16'h0000;
        rom[208][36] = 16'hFFFC;
        rom[208][37] = 16'hFFC7;
        rom[208][38] = 16'h0002;
        rom[208][39] = 16'h0005;
        rom[208][40] = 16'h002E;
        rom[208][41] = 16'h0020;
        rom[208][42] = 16'h0022;
        rom[208][43] = 16'hFFE5;
        rom[208][44] = 16'h0011;
        rom[208][45] = 16'h001F;
        rom[208][46] = 16'hFFE6;
        rom[208][47] = 16'h000E;
        rom[208][48] = 16'h0021;
        rom[208][49] = 16'h0003;
        rom[208][50] = 16'h0029;
        rom[208][51] = 16'hFFFE;
        rom[208][52] = 16'hFFCD;
        rom[208][53] = 16'h0010;
        rom[208][54] = 16'h0023;
        rom[208][55] = 16'h0005;
        rom[208][56] = 16'hFFF4;
        rom[208][57] = 16'h0000;
        rom[208][58] = 16'hFFEB;
        rom[208][59] = 16'hFFDF;
        rom[208][60] = 16'hFFC2;
        rom[208][61] = 16'hFFEF;
        rom[208][62] = 16'h001A;
        rom[208][63] = 16'h000B;
        rom[208][64] = 16'hFFD4;
        rom[208][65] = 16'hFFE8;
        rom[208][66] = 16'hFFEF;
        rom[208][67] = 16'hFFE2;
        rom[208][68] = 16'hFFD8;
        rom[208][69] = 16'hFFB3;
        rom[208][70] = 16'h000B;
        rom[208][71] = 16'hFFF8;
        rom[208][72] = 16'hFFDE;
        rom[208][73] = 16'hFFF5;
        rom[208][74] = 16'hFFEC;
        rom[208][75] = 16'hFFDB;
        rom[208][76] = 16'hFFEA;
        rom[208][77] = 16'hFFCE;
        rom[208][78] = 16'hFFEC;
        rom[208][79] = 16'hFFA3;
        rom[208][80] = 16'h0008;
        rom[208][81] = 16'hFFF9;
        rom[208][82] = 16'h0017;
        rom[208][83] = 16'h000E;
        rom[208][84] = 16'hFFA6;
        rom[208][85] = 16'h0019;
        rom[208][86] = 16'h0001;
        rom[208][87] = 16'hFFEF;
        rom[208][88] = 16'hFFF9;
        rom[208][89] = 16'h0015;
        rom[208][90] = 16'h0002;
        rom[208][91] = 16'h001F;
        rom[208][92] = 16'h0007;
        rom[208][93] = 16'h0005;
        rom[208][94] = 16'hFFDB;
        rom[208][95] = 16'h000F;
        rom[208][96] = 16'hFFFA;
        rom[208][97] = 16'h000F;
        rom[208][98] = 16'hFFD1;
        rom[208][99] = 16'hFFE6;
        rom[208][100] = 16'h0031;
        rom[208][101] = 16'h0012;
        rom[208][102] = 16'h001C;
        rom[208][103] = 16'h0013;
        rom[208][104] = 16'hFFF2;
        rom[208][105] = 16'h002E;
        rom[208][106] = 16'hFFEA;
        rom[208][107] = 16'hFFF3;
        rom[208][108] = 16'h001C;
        rom[208][109] = 16'hFFF4;
        rom[208][110] = 16'h0020;
        rom[208][111] = 16'hFFCE;
        rom[208][112] = 16'hFFE4;
        rom[208][113] = 16'hFFDE;
        rom[208][114] = 16'hFFF8;
        rom[208][115] = 16'h0016;
        rom[208][116] = 16'hFFCA;
        rom[208][117] = 16'hFFFE;
        rom[208][118] = 16'hFFEE;
        rom[208][119] = 16'h000A;
        rom[208][120] = 16'hFFE9;
        rom[208][121] = 16'h0019;
        rom[208][122] = 16'hFFF2;
        rom[208][123] = 16'hFFEB;
        rom[208][124] = 16'hFFEE;
        rom[208][125] = 16'hFFE3;
        rom[208][126] = 16'h0003;
        rom[208][127] = 16'hFFF6;
        rom[209][0] = 16'hFFEC;
        rom[209][1] = 16'h0040;
        rom[209][2] = 16'hFFD1;
        rom[209][3] = 16'hFFD3;
        rom[209][4] = 16'hFFB7;
        rom[209][5] = 16'h001B;
        rom[209][6] = 16'hFFFF;
        rom[209][7] = 16'h0024;
        rom[209][8] = 16'h0012;
        rom[209][9] = 16'hFFF7;
        rom[209][10] = 16'hFFEF;
        rom[209][11] = 16'hFFC4;
        rom[209][12] = 16'hFFE5;
        rom[209][13] = 16'hFFEE;
        rom[209][14] = 16'hFFD9;
        rom[209][15] = 16'h0007;
        rom[209][16] = 16'h0012;
        rom[209][17] = 16'h0014;
        rom[209][18] = 16'h0007;
        rom[209][19] = 16'h001F;
        rom[209][20] = 16'hFFCA;
        rom[209][21] = 16'h000B;
        rom[209][22] = 16'hFFD3;
        rom[209][23] = 16'h001D;
        rom[209][24] = 16'h0007;
        rom[209][25] = 16'h000C;
        rom[209][26] = 16'hFFDC;
        rom[209][27] = 16'hFFB5;
        rom[209][28] = 16'hFFF9;
        rom[209][29] = 16'h0005;
        rom[209][30] = 16'hFFEC;
        rom[209][31] = 16'hFFEB;
        rom[209][32] = 16'hFFD2;
        rom[209][33] = 16'h0032;
        rom[209][34] = 16'hFFED;
        rom[209][35] = 16'hFFD4;
        rom[209][36] = 16'hFFF4;
        rom[209][37] = 16'h001C;
        rom[209][38] = 16'h0006;
        rom[209][39] = 16'h001A;
        rom[209][40] = 16'h0016;
        rom[209][41] = 16'h0003;
        rom[209][42] = 16'hFFEF;
        rom[209][43] = 16'hFFC9;
        rom[209][44] = 16'hFFEB;
        rom[209][45] = 16'hFFD8;
        rom[209][46] = 16'h0012;
        rom[209][47] = 16'hFFE1;
        rom[209][48] = 16'h0002;
        rom[209][49] = 16'h0011;
        rom[209][50] = 16'hFFDC;
        rom[209][51] = 16'hFFE7;
        rom[209][52] = 16'hFFD1;
        rom[209][53] = 16'hFFE0;
        rom[209][54] = 16'hFFD6;
        rom[209][55] = 16'hFFE1;
        rom[209][56] = 16'hFFEA;
        rom[209][57] = 16'h0007;
        rom[209][58] = 16'hFFE7;
        rom[209][59] = 16'hFFF4;
        rom[209][60] = 16'h0007;
        rom[209][61] = 16'hFFD6;
        rom[209][62] = 16'h0016;
        rom[209][63] = 16'h002E;
        rom[209][64] = 16'h0010;
        rom[209][65] = 16'h0003;
        rom[209][66] = 16'hFFE0;
        rom[209][67] = 16'h0011;
        rom[209][68] = 16'h005A;
        rom[209][69] = 16'hFFFF;
        rom[209][70] = 16'hFFDC;
        rom[209][71] = 16'hFFDC;
        rom[209][72] = 16'hFFE0;
        rom[209][73] = 16'h0001;
        rom[209][74] = 16'h0021;
        rom[209][75] = 16'h0007;
        rom[209][76] = 16'hFFE7;
        rom[209][77] = 16'hFFD9;
        rom[209][78] = 16'hFFFB;
        rom[209][79] = 16'h0015;
        rom[209][80] = 16'h0021;
        rom[209][81] = 16'hFFFE;
        rom[209][82] = 16'h0019;
        rom[209][83] = 16'hFFF9;
        rom[209][84] = 16'hFFF9;
        rom[209][85] = 16'hFFFE;
        rom[209][86] = 16'h0044;
        rom[209][87] = 16'hFFF1;
        rom[209][88] = 16'h0007;
        rom[209][89] = 16'hFFE5;
        rom[209][90] = 16'h001E;
        rom[209][91] = 16'h0007;
        rom[209][92] = 16'hFFEB;
        rom[209][93] = 16'hFFF7;
        rom[209][94] = 16'h000C;
        rom[209][95] = 16'h0017;
        rom[209][96] = 16'hFFFC;
        rom[209][97] = 16'h0022;
        rom[209][98] = 16'h000E;
        rom[209][99] = 16'h0000;
        rom[209][100] = 16'h001C;
        rom[209][101] = 16'hFFF0;
        rom[209][102] = 16'hFFF5;
        rom[209][103] = 16'hFFFE;
        rom[209][104] = 16'hFFFD;
        rom[209][105] = 16'hFFEB;
        rom[209][106] = 16'hFFFF;
        rom[209][107] = 16'hFFE1;
        rom[209][108] = 16'h0016;
        rom[209][109] = 16'h0006;
        rom[209][110] = 16'hFFEA;
        rom[209][111] = 16'h000D;
        rom[209][112] = 16'hFFF2;
        rom[209][113] = 16'h0016;
        rom[209][114] = 16'hFFFE;
        rom[209][115] = 16'hFFEF;
        rom[209][116] = 16'h000C;
        rom[209][117] = 16'h0020;
        rom[209][118] = 16'hFFF7;
        rom[209][119] = 16'h0004;
        rom[209][120] = 16'hFFC7;
        rom[209][121] = 16'h0011;
        rom[209][122] = 16'hFFDA;
        rom[209][123] = 16'hFFE2;
        rom[209][124] = 16'h000C;
        rom[209][125] = 16'hFFD9;
        rom[209][126] = 16'hFFED;
        rom[209][127] = 16'hFFE1;
        rom[210][0] = 16'h000A;
        rom[210][1] = 16'h0012;
        rom[210][2] = 16'h0025;
        rom[210][3] = 16'hFFC9;
        rom[210][4] = 16'h0025;
        rom[210][5] = 16'h001D;
        rom[210][6] = 16'h0004;
        rom[210][7] = 16'hFFE4;
        rom[210][8] = 16'hFFF3;
        rom[210][9] = 16'h0010;
        rom[210][10] = 16'h000A;
        rom[210][11] = 16'h0022;
        rom[210][12] = 16'hFFE8;
        rom[210][13] = 16'hFFE5;
        rom[210][14] = 16'h0026;
        rom[210][15] = 16'h0005;
        rom[210][16] = 16'hFFEF;
        rom[210][17] = 16'hFFCA;
        rom[210][18] = 16'hFFE6;
        rom[210][19] = 16'hFFCB;
        rom[210][20] = 16'h000D;
        rom[210][21] = 16'h0020;
        rom[210][22] = 16'hFFF4;
        rom[210][23] = 16'h000B;
        rom[210][24] = 16'hFFF2;
        rom[210][25] = 16'h000F;
        rom[210][26] = 16'h0007;
        rom[210][27] = 16'h001F;
        rom[210][28] = 16'hFFDE;
        rom[210][29] = 16'hFFF1;
        rom[210][30] = 16'h000E;
        rom[210][31] = 16'hFFF4;
        rom[210][32] = 16'hFFB3;
        rom[210][33] = 16'hFFFE;
        rom[210][34] = 16'h001E;
        rom[210][35] = 16'hFFFE;
        rom[210][36] = 16'h000D;
        rom[210][37] = 16'h0002;
        rom[210][38] = 16'hFFF9;
        rom[210][39] = 16'hFFC5;
        rom[210][40] = 16'hFFEF;
        rom[210][41] = 16'h0002;
        rom[210][42] = 16'hFFEE;
        rom[210][43] = 16'hFFC4;
        rom[210][44] = 16'hFFE4;
        rom[210][45] = 16'hFFFF;
        rom[210][46] = 16'hFFFA;
        rom[210][47] = 16'hFFDE;
        rom[210][48] = 16'h0018;
        rom[210][49] = 16'h001B;
        rom[210][50] = 16'h0011;
        rom[210][51] = 16'h0010;
        rom[210][52] = 16'h0024;
        rom[210][53] = 16'hFFA6;
        rom[210][54] = 16'h005E;
        rom[210][55] = 16'hFFDD;
        rom[210][56] = 16'h0000;
        rom[210][57] = 16'hFFE5;
        rom[210][58] = 16'hFFDA;
        rom[210][59] = 16'hFFF9;
        rom[210][60] = 16'h002A;
        rom[210][61] = 16'hFFD7;
        rom[210][62] = 16'hFFE5;
        rom[210][63] = 16'hFFF1;
        rom[210][64] = 16'h0007;
        rom[210][65] = 16'hFFFE;
        rom[210][66] = 16'h002E;
        rom[210][67] = 16'hFFEB;
        rom[210][68] = 16'h0013;
        rom[210][69] = 16'hFFF9;
        rom[210][70] = 16'h0023;
        rom[210][71] = 16'h0011;
        rom[210][72] = 16'hFFE6;
        rom[210][73] = 16'h0009;
        rom[210][74] = 16'hFFEB;
        rom[210][75] = 16'h003B;
        rom[210][76] = 16'h001E;
        rom[210][77] = 16'h0003;
        rom[210][78] = 16'hFFCD;
        rom[210][79] = 16'hFFE4;
        rom[210][80] = 16'h0015;
        rom[210][81] = 16'h0011;
        rom[210][82] = 16'hFFF4;
        rom[210][83] = 16'hFFDB;
        rom[210][84] = 16'h0007;
        rom[210][85] = 16'hFFD7;
        rom[210][86] = 16'hFFD2;
        rom[210][87] = 16'h0010;
        rom[210][88] = 16'h0006;
        rom[210][89] = 16'hFFBF;
        rom[210][90] = 16'hFFF3;
        rom[210][91] = 16'h001E;
        rom[210][92] = 16'h0012;
        rom[210][93] = 16'hFFF0;
        rom[210][94] = 16'hFFD4;
        rom[210][95] = 16'hFFD1;
        rom[210][96] = 16'hFFC8;
        rom[210][97] = 16'hFFFB;
        rom[210][98] = 16'h001A;
        rom[210][99] = 16'h0019;
        rom[210][100] = 16'hFFFB;
        rom[210][101] = 16'h0011;
        rom[210][102] = 16'h0019;
        rom[210][103] = 16'h002D;
        rom[210][104] = 16'h000A;
        rom[210][105] = 16'h0001;
        rom[210][106] = 16'h001B;
        rom[210][107] = 16'h0029;
        rom[210][108] = 16'hFFF1;
        rom[210][109] = 16'hFFD3;
        rom[210][110] = 16'hFFFE;
        rom[210][111] = 16'h0002;
        rom[210][112] = 16'hFFFC;
        rom[210][113] = 16'hFFF1;
        rom[210][114] = 16'h0036;
        rom[210][115] = 16'hFFF2;
        rom[210][116] = 16'h0007;
        rom[210][117] = 16'h0018;
        rom[210][118] = 16'hFFE9;
        rom[210][119] = 16'h0031;
        rom[210][120] = 16'hFFEE;
        rom[210][121] = 16'hFFEA;
        rom[210][122] = 16'h0014;
        rom[210][123] = 16'h0012;
        rom[210][124] = 16'hFFDA;
        rom[210][125] = 16'hFFF9;
        rom[210][126] = 16'hFFEC;
        rom[210][127] = 16'hFFF7;
        rom[211][0] = 16'hFFFB;
        rom[211][1] = 16'h000F;
        rom[211][2] = 16'hFFFF;
        rom[211][3] = 16'h0002;
        rom[211][4] = 16'hFFFD;
        rom[211][5] = 16'hFFED;
        rom[211][6] = 16'hFFE0;
        rom[211][7] = 16'h000F;
        rom[211][8] = 16'hFFC6;
        rom[211][9] = 16'hFFE7;
        rom[211][10] = 16'hFFE3;
        rom[211][11] = 16'hFFEF;
        rom[211][12] = 16'hFFFE;
        rom[211][13] = 16'hFFF6;
        rom[211][14] = 16'h0004;
        rom[211][15] = 16'hFFFC;
        rom[211][16] = 16'hFFD6;
        rom[211][17] = 16'h0019;
        rom[211][18] = 16'hFFEE;
        rom[211][19] = 16'h0024;
        rom[211][20] = 16'hFFF9;
        rom[211][21] = 16'h0016;
        rom[211][22] = 16'hFFEA;
        rom[211][23] = 16'h001C;
        rom[211][24] = 16'hFFFF;
        rom[211][25] = 16'hFFFA;
        rom[211][26] = 16'hFFEA;
        rom[211][27] = 16'h0005;
        rom[211][28] = 16'h0048;
        rom[211][29] = 16'h0011;
        rom[211][30] = 16'hFFFF;
        rom[211][31] = 16'hFFF8;
        rom[211][32] = 16'hFFF8;
        rom[211][33] = 16'hFFFA;
        rom[211][34] = 16'hFFE9;
        rom[211][35] = 16'hFFE6;
        rom[211][36] = 16'hFFED;
        rom[211][37] = 16'h0010;
        rom[211][38] = 16'hFFE9;
        rom[211][39] = 16'hFFDB;
        rom[211][40] = 16'h0011;
        rom[211][41] = 16'h000C;
        rom[211][42] = 16'h0010;
        rom[211][43] = 16'hFFE0;
        rom[211][44] = 16'hFFDC;
        rom[211][45] = 16'hFFEE;
        rom[211][46] = 16'hFFFB;
        rom[211][47] = 16'hFFF4;
        rom[211][48] = 16'hFFBA;
        rom[211][49] = 16'hFFE5;
        rom[211][50] = 16'hFFDA;
        rom[211][51] = 16'hFFD7;
        rom[211][52] = 16'h001C;
        rom[211][53] = 16'h0011;
        rom[211][54] = 16'h0003;
        rom[211][55] = 16'h0042;
        rom[211][56] = 16'h001C;
        rom[211][57] = 16'hFFD9;
        rom[211][58] = 16'hFFD1;
        rom[211][59] = 16'h0011;
        rom[211][60] = 16'hFFF5;
        rom[211][61] = 16'h0015;
        rom[211][62] = 16'hFFF5;
        rom[211][63] = 16'hFFD4;
        rom[211][64] = 16'h0007;
        rom[211][65] = 16'hFFEA;
        rom[211][66] = 16'hFFFE;
        rom[211][67] = 16'h001C;
        rom[211][68] = 16'hFFFA;
        rom[211][69] = 16'hFFF4;
        rom[211][70] = 16'hFFEF;
        rom[211][71] = 16'hFFD7;
        rom[211][72] = 16'hFFF9;
        rom[211][73] = 16'h0010;
        rom[211][74] = 16'hFFE0;
        rom[211][75] = 16'h000F;
        rom[211][76] = 16'h001D;
        rom[211][77] = 16'h000F;
        rom[211][78] = 16'hFFD9;
        rom[211][79] = 16'hFFE0;
        rom[211][80] = 16'h000C;
        rom[211][81] = 16'hFFE9;
        rom[211][82] = 16'h002E;
        rom[211][83] = 16'h001E;
        rom[211][84] = 16'hFFE4;
        rom[211][85] = 16'h0009;
        rom[211][86] = 16'hFFFE;
        rom[211][87] = 16'hFFF2;
        rom[211][88] = 16'hFFC8;
        rom[211][89] = 16'h000B;
        rom[211][90] = 16'h001C;
        rom[211][91] = 16'hFFB0;
        rom[211][92] = 16'h000F;
        rom[211][93] = 16'hFFF2;
        rom[211][94] = 16'h0003;
        rom[211][95] = 16'h001B;
        rom[211][96] = 16'hFFC6;
        rom[211][97] = 16'hFFD7;
        rom[211][98] = 16'hFFE7;
        rom[211][99] = 16'hFFEC;
        rom[211][100] = 16'hFFFC;
        rom[211][101] = 16'h001F;
        rom[211][102] = 16'hFFDE;
        rom[211][103] = 16'hFFF9;
        rom[211][104] = 16'h0004;
        rom[211][105] = 16'hFFF7;
        rom[211][106] = 16'h0026;
        rom[211][107] = 16'hFFF4;
        rom[211][108] = 16'hFFD9;
        rom[211][109] = 16'hFFFD;
        rom[211][110] = 16'h0010;
        rom[211][111] = 16'h0016;
        rom[211][112] = 16'h001D;
        rom[211][113] = 16'hFFF0;
        rom[211][114] = 16'hFFEF;
        rom[211][115] = 16'hFFF1;
        rom[211][116] = 16'hFFF6;
        rom[211][117] = 16'h001A;
        rom[211][118] = 16'h0033;
        rom[211][119] = 16'hFFFE;
        rom[211][120] = 16'h0007;
        rom[211][121] = 16'hFFF6;
        rom[211][122] = 16'h0009;
        rom[211][123] = 16'h0009;
        rom[211][124] = 16'hFFF4;
        rom[211][125] = 16'hFFE5;
        rom[211][126] = 16'h001B;
        rom[211][127] = 16'hFFCF;
        rom[212][0] = 16'h001B;
        rom[212][1] = 16'hFFD7;
        rom[212][2] = 16'hFFEF;
        rom[212][3] = 16'hFFF4;
        rom[212][4] = 16'hFFE1;
        rom[212][5] = 16'hFFE4;
        rom[212][6] = 16'hFFE5;
        rom[212][7] = 16'h003D;
        rom[212][8] = 16'hFFFC;
        rom[212][9] = 16'h0013;
        rom[212][10] = 16'h002A;
        rom[212][11] = 16'h0024;
        rom[212][12] = 16'h0006;
        rom[212][13] = 16'h0030;
        rom[212][14] = 16'hFFEF;
        rom[212][15] = 16'hFFEA;
        rom[212][16] = 16'hFF98;
        rom[212][17] = 16'h0011;
        rom[212][18] = 16'h000C;
        rom[212][19] = 16'hFFEA;
        rom[212][20] = 16'hFFE4;
        rom[212][21] = 16'h0026;
        rom[212][22] = 16'h0003;
        rom[212][23] = 16'h0009;
        rom[212][24] = 16'h0007;
        rom[212][25] = 16'hFFF2;
        rom[212][26] = 16'hFFE7;
        rom[212][27] = 16'hFFC5;
        rom[212][28] = 16'h000B;
        rom[212][29] = 16'h001B;
        rom[212][30] = 16'h0011;
        rom[212][31] = 16'h0019;
        rom[212][32] = 16'h0004;
        rom[212][33] = 16'h001D;
        rom[212][34] = 16'hFFE0;
        rom[212][35] = 16'h0005;
        rom[212][36] = 16'h0003;
        rom[212][37] = 16'hFFF4;
        rom[212][38] = 16'h0007;
        rom[212][39] = 16'h0030;
        rom[212][40] = 16'h0016;
        rom[212][41] = 16'h001B;
        rom[212][42] = 16'hFFEB;
        rom[212][43] = 16'h000C;
        rom[212][44] = 16'h0011;
        rom[212][45] = 16'hFFFB;
        rom[212][46] = 16'hFFE7;
        rom[212][47] = 16'hFFEC;
        rom[212][48] = 16'hFFC7;
        rom[212][49] = 16'hFFAE;
        rom[212][50] = 16'hFFE4;
        rom[212][51] = 16'h0018;
        rom[212][52] = 16'h0007;
        rom[212][53] = 16'hFFFE;
        rom[212][54] = 16'hFFE3;
        rom[212][55] = 16'hFFD3;
        rom[212][56] = 16'hFFFF;
        rom[212][57] = 16'h0001;
        rom[212][58] = 16'h0019;
        rom[212][59] = 16'hFFE1;
        rom[212][60] = 16'hFFAD;
        rom[212][61] = 16'h0002;
        rom[212][62] = 16'hFFDE;
        rom[212][63] = 16'h000C;
        rom[212][64] = 16'hFFF5;
        rom[212][65] = 16'hFFFA;
        rom[212][66] = 16'hFFE4;
        rom[212][67] = 16'hFFD0;
        rom[212][68] = 16'hFFF3;
        rom[212][69] = 16'hFFA8;
        rom[212][70] = 16'hFFFF;
        rom[212][71] = 16'hFFF9;
        rom[212][72] = 16'h0012;
        rom[212][73] = 16'hFFCA;
        rom[212][74] = 16'h0031;
        rom[212][75] = 16'h0011;
        rom[212][76] = 16'h0015;
        rom[212][77] = 16'h0021;
        rom[212][78] = 16'h0013;
        rom[212][79] = 16'hFFE6;
        rom[212][80] = 16'h0000;
        rom[212][81] = 16'hFFDC;
        rom[212][82] = 16'hFFDE;
        rom[212][83] = 16'h0007;
        rom[212][84] = 16'hFFC1;
        rom[212][85] = 16'hFFF5;
        rom[212][86] = 16'h003E;
        rom[212][87] = 16'hFFD1;
        rom[212][88] = 16'hFFF5;
        rom[212][89] = 16'hFFFA;
        rom[212][90] = 16'hFFE0;
        rom[212][91] = 16'hFFB0;
        rom[212][92] = 16'hFFC0;
        rom[212][93] = 16'hFFD1;
        rom[212][94] = 16'h000B;
        rom[212][95] = 16'hFFDC;
        rom[212][96] = 16'h0014;
        rom[212][97] = 16'h000C;
        rom[212][98] = 16'hFF9B;
        rom[212][99] = 16'hFFD2;
        rom[212][100] = 16'h001B;
        rom[212][101] = 16'hFFF7;
        rom[212][102] = 16'hFFF1;
        rom[212][103] = 16'h000A;
        rom[212][104] = 16'hFFF7;
        rom[212][105] = 16'hFFEA;
        rom[212][106] = 16'h0011;
        rom[212][107] = 16'hFFFD;
        rom[212][108] = 16'hFFEF;
        rom[212][109] = 16'h0006;
        rom[212][110] = 16'hFFD0;
        rom[212][111] = 16'hFFC4;
        rom[212][112] = 16'h000A;
        rom[212][113] = 16'hFFF9;
        rom[212][114] = 16'hFFD3;
        rom[212][115] = 16'hFFF8;
        rom[212][116] = 16'hFFFE;
        rom[212][117] = 16'hFFF9;
        rom[212][118] = 16'h0013;
        rom[212][119] = 16'hFFF8;
        rom[212][120] = 16'hFFF0;
        rom[212][121] = 16'h0011;
        rom[212][122] = 16'hFFF2;
        rom[212][123] = 16'hFFC7;
        rom[212][124] = 16'hFFD8;
        rom[212][125] = 16'h000C;
        rom[212][126] = 16'h0007;
        rom[212][127] = 16'hFFE4;
        rom[213][0] = 16'hFFDF;
        rom[213][1] = 16'hFFFE;
        rom[213][2] = 16'h0012;
        rom[213][3] = 16'hFFF4;
        rom[213][4] = 16'hFFF3;
        rom[213][5] = 16'hFFEF;
        rom[213][6] = 16'hFFEF;
        rom[213][7] = 16'hFFE1;
        rom[213][8] = 16'hFFEF;
        rom[213][9] = 16'h0007;
        rom[213][10] = 16'hFFCE;
        rom[213][11] = 16'h000B;
        rom[213][12] = 16'hFFE3;
        rom[213][13] = 16'h0001;
        rom[213][14] = 16'hFFF6;
        rom[213][15] = 16'h0016;
        rom[213][16] = 16'h001D;
        rom[213][17] = 16'h0007;
        rom[213][18] = 16'hFFEB;
        rom[213][19] = 16'hFFED;
        rom[213][20] = 16'hFFDC;
        rom[213][21] = 16'hFFF9;
        rom[213][22] = 16'hFFEF;
        rom[213][23] = 16'hFFA3;
        rom[213][24] = 16'h002B;
        rom[213][25] = 16'hFFBA;
        rom[213][26] = 16'hFFE5;
        rom[213][27] = 16'hFFDE;
        rom[213][28] = 16'hFFF1;
        rom[213][29] = 16'h0000;
        rom[213][30] = 16'hFFE6;
        rom[213][31] = 16'h000B;
        rom[213][32] = 16'h0007;
        rom[213][33] = 16'hFFB1;
        rom[213][34] = 16'hFFE6;
        rom[213][35] = 16'h0034;
        rom[213][36] = 16'hFFE4;
        rom[213][37] = 16'hFFF3;
        rom[213][38] = 16'hFFF1;
        rom[213][39] = 16'hFFFD;
        rom[213][40] = 16'h0018;
        rom[213][41] = 16'h0016;
        rom[213][42] = 16'hFFAD;
        rom[213][43] = 16'h0028;
        rom[213][44] = 16'h000A;
        rom[213][45] = 16'hFFF9;
        rom[213][46] = 16'hFFF4;
        rom[213][47] = 16'hFFF6;
        rom[213][48] = 16'h000C;
        rom[213][49] = 16'h0002;
        rom[213][50] = 16'hFFE1;
        rom[213][51] = 16'h0016;
        rom[213][52] = 16'hFFFC;
        rom[213][53] = 16'h0016;
        rom[213][54] = 16'h0016;
        rom[213][55] = 16'hFFD4;
        rom[213][56] = 16'h001D;
        rom[213][57] = 16'hFFDA;
        rom[213][58] = 16'h000F;
        rom[213][59] = 16'hFFCA;
        rom[213][60] = 16'h001C;
        rom[213][61] = 16'hFFF7;
        rom[213][62] = 16'hFFF3;
        rom[213][63] = 16'hFFD4;
        rom[213][64] = 16'hFFEA;
        rom[213][65] = 16'hFFFE;
        rom[213][66] = 16'hFFDC;
        rom[213][67] = 16'hFFEF;
        rom[213][68] = 16'h0023;
        rom[213][69] = 16'hFFD4;
        rom[213][70] = 16'h0019;
        rom[213][71] = 16'h001E;
        rom[213][72] = 16'hFFFC;
        rom[213][73] = 16'hFFFB;
        rom[213][74] = 16'h0007;
        rom[213][75] = 16'hFFEA;
        rom[213][76] = 16'h0003;
        rom[213][77] = 16'h0003;
        rom[213][78] = 16'h0026;
        rom[213][79] = 16'hFFEA;
        rom[213][80] = 16'h001F;
        rom[213][81] = 16'h0002;
        rom[213][82] = 16'hFF9A;
        rom[213][83] = 16'hFFF2;
        rom[213][84] = 16'h0002;
        rom[213][85] = 16'h0012;
        rom[213][86] = 16'hFFF5;
        rom[213][87] = 16'hFFFF;
        rom[213][88] = 16'hFFE7;
        rom[213][89] = 16'h0000;
        rom[213][90] = 16'hFFB4;
        rom[213][91] = 16'hFFFE;
        rom[213][92] = 16'h000E;
        rom[213][93] = 16'hFFCC;
        rom[213][94] = 16'h000F;
        rom[213][95] = 16'hFFE4;
        rom[213][96] = 16'h0032;
        rom[213][97] = 16'hFFDD;
        rom[213][98] = 16'hFFEF;
        rom[213][99] = 16'h0004;
        rom[213][100] = 16'hFFDB;
        rom[213][101] = 16'hFFE5;
        rom[213][102] = 16'hFFD4;
        rom[213][103] = 16'hFFAF;
        rom[213][104] = 16'hFFE2;
        rom[213][105] = 16'hFFC4;
        rom[213][106] = 16'hFFF4;
        rom[213][107] = 16'hFFEC;
        rom[213][108] = 16'h000D;
        rom[213][109] = 16'h000C;
        rom[213][110] = 16'hFFD2;
        rom[213][111] = 16'h0014;
        rom[213][112] = 16'h0002;
        rom[213][113] = 16'hFFD2;
        rom[213][114] = 16'hFFE1;
        rom[213][115] = 16'hFFEA;
        rom[213][116] = 16'hFFCE;
        rom[213][117] = 16'h0005;
        rom[213][118] = 16'h0003;
        rom[213][119] = 16'h0017;
        rom[213][120] = 16'h000B;
        rom[213][121] = 16'hFFBF;
        rom[213][122] = 16'h001B;
        rom[213][123] = 16'hFFE4;
        rom[213][124] = 16'h002F;
        rom[213][125] = 16'hFFF8;
        rom[213][126] = 16'h0003;
        rom[213][127] = 16'hFFEF;
        rom[214][0] = 16'h002B;
        rom[214][1] = 16'hFFB1;
        rom[214][2] = 16'h0018;
        rom[214][3] = 16'h0013;
        rom[214][4] = 16'hFFD1;
        rom[214][5] = 16'hFFF6;
        rom[214][6] = 16'h000B;
        rom[214][7] = 16'h0018;
        rom[214][8] = 16'hFFFF;
        rom[214][9] = 16'hFFEC;
        rom[214][10] = 16'hFFE1;
        rom[214][11] = 16'h001F;
        rom[214][12] = 16'hFFF9;
        rom[214][13] = 16'h0014;
        rom[214][14] = 16'hFFCA;
        rom[214][15] = 16'hFFF3;
        rom[214][16] = 16'h0016;
        rom[214][17] = 16'h0007;
        rom[214][18] = 16'h001B;
        rom[214][19] = 16'hFFBD;
        rom[214][20] = 16'h0032;
        rom[214][21] = 16'hFFD3;
        rom[214][22] = 16'hFFD7;
        rom[214][23] = 16'h0015;
        rom[214][24] = 16'h0011;
        rom[214][25] = 16'h001A;
        rom[214][26] = 16'h0007;
        rom[214][27] = 16'hFFD6;
        rom[214][28] = 16'hFFAF;
        rom[214][29] = 16'hFFCF;
        rom[214][30] = 16'hFFF6;
        rom[214][31] = 16'h0024;
        rom[214][32] = 16'h0028;
        rom[214][33] = 16'hFFD2;
        rom[214][34] = 16'h002D;
        rom[214][35] = 16'h0010;
        rom[214][36] = 16'h0020;
        rom[214][37] = 16'hFFDD;
        rom[214][38] = 16'h0004;
        rom[214][39] = 16'hFFEB;
        rom[214][40] = 16'hFFE6;
        rom[214][41] = 16'hFFE5;
        rom[214][42] = 16'hFFF1;
        rom[214][43] = 16'hFFE1;
        rom[214][44] = 16'h0020;
        rom[214][45] = 16'h000C;
        rom[214][46] = 16'hFFE6;
        rom[214][47] = 16'hFFD9;
        rom[214][48] = 16'h001F;
        rom[214][49] = 16'h001B;
        rom[214][50] = 16'h0029;
        rom[214][51] = 16'h0030;
        rom[214][52] = 16'hFFEB;
        rom[214][53] = 16'h0002;
        rom[214][54] = 16'hFFEB;
        rom[214][55] = 16'h0004;
        rom[214][56] = 16'hFFEF;
        rom[214][57] = 16'h0052;
        rom[214][58] = 16'hFFC8;
        rom[214][59] = 16'h001B;
        rom[214][60] = 16'hFFF1;
        rom[214][61] = 16'hFFF7;
        rom[214][62] = 16'hFFD2;
        rom[214][63] = 16'h0032;
        rom[214][64] = 16'h0007;
        rom[214][65] = 16'hFFC7;
        rom[214][66] = 16'hFFF1;
        rom[214][67] = 16'hFFB0;
        rom[214][68] = 16'hFFEA;
        rom[214][69] = 16'hFFCD;
        rom[214][70] = 16'hFFED;
        rom[214][71] = 16'h0014;
        rom[214][72] = 16'h0016;
        rom[214][73] = 16'hFFAD;
        rom[214][74] = 16'h001F;
        rom[214][75] = 16'hFFC2;
        rom[214][76] = 16'h0024;
        rom[214][77] = 16'hFFB5;
        rom[214][78] = 16'hFFFF;
        rom[214][79] = 16'hFFC4;
        rom[214][80] = 16'hFFE9;
        rom[214][81] = 16'hFFFE;
        rom[214][82] = 16'hFFEB;
        rom[214][83] = 16'h0014;
        rom[214][84] = 16'h0002;
        rom[214][85] = 16'h002D;
        rom[214][86] = 16'hFFFE;
        rom[214][87] = 16'h0016;
        rom[214][88] = 16'h003A;
        rom[214][89] = 16'hFFF0;
        rom[214][90] = 16'hFFE6;
        rom[214][91] = 16'hFFE6;
        rom[214][92] = 16'hFFE4;
        rom[214][93] = 16'hFFD8;
        rom[214][94] = 16'hFFF1;
        rom[214][95] = 16'hFFD6;
        rom[214][96] = 16'h0007;
        rom[214][97] = 16'h0009;
        rom[214][98] = 16'hFFC4;
        rom[214][99] = 16'h0007;
        rom[214][100] = 16'hFFD1;
        rom[214][101] = 16'hFFEF;
        rom[214][102] = 16'h001A;
        rom[214][103] = 16'h0018;
        rom[214][104] = 16'hFFE2;
        rom[214][105] = 16'hFFD8;
        rom[214][106] = 16'hFFE3;
        rom[214][107] = 16'h0010;
        rom[214][108] = 16'hFFF8;
        rom[214][109] = 16'h000E;
        rom[214][110] = 16'hFFE5;
        rom[214][111] = 16'hFFD8;
        rom[214][112] = 16'hFFE8;
        rom[214][113] = 16'h001F;
        rom[214][114] = 16'h0010;
        rom[214][115] = 16'h0002;
        rom[214][116] = 16'hFFF0;
        rom[214][117] = 16'hFFE7;
        rom[214][118] = 16'hFFEB;
        rom[214][119] = 16'hFFEF;
        rom[214][120] = 16'h0024;
        rom[214][121] = 16'hFFE1;
        rom[214][122] = 16'h001B;
        rom[214][123] = 16'h000B;
        rom[214][124] = 16'hFFE5;
        rom[214][125] = 16'hFFD7;
        rom[214][126] = 16'hFFF4;
        rom[214][127] = 16'h0001;
        rom[215][0] = 16'hFFE3;
        rom[215][1] = 16'h0016;
        rom[215][2] = 16'hFFCE;
        rom[215][3] = 16'h0016;
        rom[215][4] = 16'h0007;
        rom[215][5] = 16'h0009;
        rom[215][6] = 16'hFFF9;
        rom[215][7] = 16'hFFFE;
        rom[215][8] = 16'hFFFE;
        rom[215][9] = 16'h002C;
        rom[215][10] = 16'h0019;
        rom[215][11] = 16'h002D;
        rom[215][12] = 16'h0010;
        rom[215][13] = 16'h000F;
        rom[215][14] = 16'h0033;
        rom[215][15] = 16'hFFBC;
        rom[215][16] = 16'h0011;
        rom[215][17] = 16'hFFFC;
        rom[215][18] = 16'hFFF4;
        rom[215][19] = 16'h000C;
        rom[215][20] = 16'hFFE8;
        rom[215][21] = 16'hFFCE;
        rom[215][22] = 16'hFFFC;
        rom[215][23] = 16'h001F;
        rom[215][24] = 16'h0029;
        rom[215][25] = 16'hFFCD;
        rom[215][26] = 16'hFFEF;
        rom[215][27] = 16'hFFF3;
        rom[215][28] = 16'h0019;
        rom[215][29] = 16'h0014;
        rom[215][30] = 16'h002F;
        rom[215][31] = 16'hFFE7;
        rom[215][32] = 16'h0024;
        rom[215][33] = 16'hFFEA;
        rom[215][34] = 16'hFFD7;
        rom[215][35] = 16'h001B;
        rom[215][36] = 16'hFFFB;
        rom[215][37] = 16'hFFD7;
        rom[215][38] = 16'hFFE8;
        rom[215][39] = 16'h0012;
        rom[215][40] = 16'hFFF3;
        rom[215][41] = 16'hFFDA;
        rom[215][42] = 16'hFFF2;
        rom[215][43] = 16'hFFE8;
        rom[215][44] = 16'hFFE8;
        rom[215][45] = 16'hFFF1;
        rom[215][46] = 16'h002D;
        rom[215][47] = 16'h0010;
        rom[215][48] = 16'hFFF2;
        rom[215][49] = 16'hFFE2;
        rom[215][50] = 16'hFFFC;
        rom[215][51] = 16'hFFC0;
        rom[215][52] = 16'hFFC0;
        rom[215][53] = 16'h0004;
        rom[215][54] = 16'h0016;
        rom[215][55] = 16'hFFDF;
        rom[215][56] = 16'h0000;
        rom[215][57] = 16'hFFD5;
        rom[215][58] = 16'hFFFD;
        rom[215][59] = 16'h002E;
        rom[215][60] = 16'h000F;
        rom[215][61] = 16'h0029;
        rom[215][62] = 16'h002E;
        rom[215][63] = 16'hFFF5;
        rom[215][64] = 16'hFFFE;
        rom[215][65] = 16'hFFF8;
        rom[215][66] = 16'h0013;
        rom[215][67] = 16'hFFDE;
        rom[215][68] = 16'hFFF5;
        rom[215][69] = 16'hFFF4;
        rom[215][70] = 16'hFFEA;
        rom[215][71] = 16'hFFF3;
        rom[215][72] = 16'h0012;
        rom[215][73] = 16'h0024;
        rom[215][74] = 16'hFFCA;
        rom[215][75] = 16'hFFDE;
        rom[215][76] = 16'hFFE5;
        rom[215][77] = 16'h0035;
        rom[215][78] = 16'h002E;
        rom[215][79] = 16'h0008;
        rom[215][80] = 16'hFFFF;
        rom[215][81] = 16'hFFE2;
        rom[215][82] = 16'h0029;
        rom[215][83] = 16'h0026;
        rom[215][84] = 16'hFFF6;
        rom[215][85] = 16'h0018;
        rom[215][86] = 16'h003A;
        rom[215][87] = 16'h0010;
        rom[215][88] = 16'hFFE1;
        rom[215][89] = 16'h0005;
        rom[215][90] = 16'hFFED;
        rom[215][91] = 16'h0002;
        rom[215][92] = 16'hFFF5;
        rom[215][93] = 16'h002A;
        rom[215][94] = 16'hFFED;
        rom[215][95] = 16'h0013;
        rom[215][96] = 16'h0012;
        rom[215][97] = 16'hFFE0;
        rom[215][98] = 16'h000A;
        rom[215][99] = 16'hFFFA;
        rom[215][100] = 16'hFFFB;
        rom[215][101] = 16'hFFD7;
        rom[215][102] = 16'hFFE2;
        rom[215][103] = 16'hFFE3;
        rom[215][104] = 16'hFFBE;
        rom[215][105] = 16'hFFF8;
        rom[215][106] = 16'h0007;
        rom[215][107] = 16'hFFEF;
        rom[215][108] = 16'hFFF8;
        rom[215][109] = 16'h0015;
        rom[215][110] = 16'h0002;
        rom[215][111] = 16'h0051;
        rom[215][112] = 16'hFFD8;
        rom[215][113] = 16'hFFD7;
        rom[215][114] = 16'hFFD7;
        rom[215][115] = 16'hFFE9;
        rom[215][116] = 16'h0000;
        rom[215][117] = 16'h0003;
        rom[215][118] = 16'h0033;
        rom[215][119] = 16'hFFE4;
        rom[215][120] = 16'h001A;
        rom[215][121] = 16'h003A;
        rom[215][122] = 16'h0033;
        rom[215][123] = 16'h0002;
        rom[215][124] = 16'h000D;
        rom[215][125] = 16'hFFC3;
        rom[215][126] = 16'hFFFB;
        rom[215][127] = 16'hFFF4;
        rom[216][0] = 16'hFFED;
        rom[216][1] = 16'h0005;
        rom[216][2] = 16'h0005;
        rom[216][3] = 16'h001B;
        rom[216][4] = 16'hFFED;
        rom[216][5] = 16'h0029;
        rom[216][6] = 16'hFFD6;
        rom[216][7] = 16'hFFF7;
        rom[216][8] = 16'h0018;
        rom[216][9] = 16'hFFF3;
        rom[216][10] = 16'hFFDD;
        rom[216][11] = 16'h0004;
        rom[216][12] = 16'hFFC4;
        rom[216][13] = 16'hFFDB;
        rom[216][14] = 16'h0002;
        rom[216][15] = 16'h001B;
        rom[216][16] = 16'hFFF9;
        rom[216][17] = 16'hFFE5;
        rom[216][18] = 16'hFFFC;
        rom[216][19] = 16'hFFEF;
        rom[216][20] = 16'hFFDA;
        rom[216][21] = 16'h0037;
        rom[216][22] = 16'h0066;
        rom[216][23] = 16'h0025;
        rom[216][24] = 16'h000C;
        rom[216][25] = 16'hFFEE;
        rom[216][26] = 16'h000F;
        rom[216][27] = 16'hFFF0;
        rom[216][28] = 16'h000E;
        rom[216][29] = 16'hFFD2;
        rom[216][30] = 16'h0003;
        rom[216][31] = 16'hFFF9;
        rom[216][32] = 16'hFFD2;
        rom[216][33] = 16'hFFC8;
        rom[216][34] = 16'h0015;
        rom[216][35] = 16'h0006;
        rom[216][36] = 16'h0010;
        rom[216][37] = 16'hFFF2;
        rom[216][38] = 16'hFFF9;
        rom[216][39] = 16'h0037;
        rom[216][40] = 16'hFFBF;
        rom[216][41] = 16'h003D;
        rom[216][42] = 16'hFFB6;
        rom[216][43] = 16'h0033;
        rom[216][44] = 16'hFFEC;
        rom[216][45] = 16'h0021;
        rom[216][46] = 16'hFFF6;
        rom[216][47] = 16'h002E;
        rom[216][48] = 16'hFFE1;
        rom[216][49] = 16'hFFD6;
        rom[216][50] = 16'hFFF9;
        rom[216][51] = 16'hFFD7;
        rom[216][52] = 16'h0016;
        rom[216][53] = 16'hFFFE;
        rom[216][54] = 16'h0006;
        rom[216][55] = 16'h0029;
        rom[216][56] = 16'hFFF5;
        rom[216][57] = 16'hFFA6;
        rom[216][58] = 16'hFFEF;
        rom[216][59] = 16'hFFE3;
        rom[216][60] = 16'h001F;
        rom[216][61] = 16'h0000;
        rom[216][62] = 16'h001D;
        rom[216][63] = 16'h0005;
        rom[216][64] = 16'hFFA4;
        rom[216][65] = 16'h0008;
        rom[216][66] = 16'hFFC5;
        rom[216][67] = 16'hFFE6;
        rom[216][68] = 16'hFFD4;
        rom[216][69] = 16'h001F;
        rom[216][70] = 16'h0011;
        rom[216][71] = 16'h001B;
        rom[216][72] = 16'hFFFD;
        rom[216][73] = 16'hFFF4;
        rom[216][74] = 16'hFFEA;
        rom[216][75] = 16'h0010;
        rom[216][76] = 16'hFFE7;
        rom[216][77] = 16'hFFE3;
        rom[216][78] = 16'h0011;
        rom[216][79] = 16'hFFE0;
        rom[216][80] = 16'hFFFE;
        rom[216][81] = 16'h0003;
        rom[216][82] = 16'hFFEF;
        rom[216][83] = 16'h0019;
        rom[216][84] = 16'h0001;
        rom[216][85] = 16'hFFFB;
        rom[216][86] = 16'hFFB2;
        rom[216][87] = 16'h001F;
        rom[216][88] = 16'h0029;
        rom[216][89] = 16'h000D;
        rom[216][90] = 16'hFFFD;
        rom[216][91] = 16'h0001;
        rom[216][92] = 16'h0004;
        rom[216][93] = 16'h000F;
        rom[216][94] = 16'hFFFE;
        rom[216][95] = 16'hFFE0;
        rom[216][96] = 16'h0011;
        rom[216][97] = 16'hFFE0;
        rom[216][98] = 16'hFFF3;
        rom[216][99] = 16'h002F;
        rom[216][100] = 16'hFFDA;
        rom[216][101] = 16'hFFDC;
        rom[216][102] = 16'hFFA3;
        rom[216][103] = 16'hFFCE;
        rom[216][104] = 16'hFFD7;
        rom[216][105] = 16'hFFAB;
        rom[216][106] = 16'hFFE8;
        rom[216][107] = 16'h0019;
        rom[216][108] = 16'hFFF4;
        rom[216][109] = 16'hFFF7;
        rom[216][110] = 16'hFFEF;
        rom[216][111] = 16'h0036;
        rom[216][112] = 16'hFFFA;
        rom[216][113] = 16'h002C;
        rom[216][114] = 16'hFFF4;
        rom[216][115] = 16'h003E;
        rom[216][116] = 16'hFFF9;
        rom[216][117] = 16'hFFC9;
        rom[216][118] = 16'hFFF3;
        rom[216][119] = 16'h0021;
        rom[216][120] = 16'hFFD7;
        rom[216][121] = 16'hFFEF;
        rom[216][122] = 16'h0011;
        rom[216][123] = 16'h0002;
        rom[216][124] = 16'h001A;
        rom[216][125] = 16'hFFF8;
        rom[216][126] = 16'h0020;
        rom[216][127] = 16'h0007;
        rom[217][0] = 16'h0007;
        rom[217][1] = 16'h0006;
        rom[217][2] = 16'hFFF5;
        rom[217][3] = 16'h000C;
        rom[217][4] = 16'h0003;
        rom[217][5] = 16'h0014;
        rom[217][6] = 16'h002A;
        rom[217][7] = 16'h0007;
        rom[217][8] = 16'hFFDC;
        rom[217][9] = 16'hFFC7;
        rom[217][10] = 16'hFFD0;
        rom[217][11] = 16'h0006;
        rom[217][12] = 16'hFFC8;
        rom[217][13] = 16'hFFCB;
        rom[217][14] = 16'hFFD7;
        rom[217][15] = 16'h0011;
        rom[217][16] = 16'h0014;
        rom[217][17] = 16'hFFE7;
        rom[217][18] = 16'hFFF9;
        rom[217][19] = 16'hFFE1;
        rom[217][20] = 16'hFFD8;
        rom[217][21] = 16'hFFF4;
        rom[217][22] = 16'hFFE7;
        rom[217][23] = 16'h0010;
        rom[217][24] = 16'hFFE6;
        rom[217][25] = 16'hFFD9;
        rom[217][26] = 16'hFFE9;
        rom[217][27] = 16'hFF96;
        rom[217][28] = 16'hFFE3;
        rom[217][29] = 16'hFFBC;
        rom[217][30] = 16'hFFEE;
        rom[217][31] = 16'hFFF8;
        rom[217][32] = 16'h0000;
        rom[217][33] = 16'hFFA3;
        rom[217][34] = 16'h000A;
        rom[217][35] = 16'h0014;
        rom[217][36] = 16'h0011;
        rom[217][37] = 16'hFFE2;
        rom[217][38] = 16'hFFD9;
        rom[217][39] = 16'h0024;
        rom[217][40] = 16'hFFD4;
        rom[217][41] = 16'h0003;
        rom[217][42] = 16'hFFA9;
        rom[217][43] = 16'h0016;
        rom[217][44] = 16'hFFF6;
        rom[217][45] = 16'hFFF6;
        rom[217][46] = 16'h0035;
        rom[217][47] = 16'hFFD2;
        rom[217][48] = 16'h0020;
        rom[217][49] = 16'h0019;
        rom[217][50] = 16'h0024;
        rom[217][51] = 16'hFFEC;
        rom[217][52] = 16'h0010;
        rom[217][53] = 16'h0011;
        rom[217][54] = 16'h0015;
        rom[217][55] = 16'hFFF2;
        rom[217][56] = 16'hFFEA;
        rom[217][57] = 16'h0016;
        rom[217][58] = 16'hFFEF;
        rom[217][59] = 16'hFFB3;
        rom[217][60] = 16'h000D;
        rom[217][61] = 16'hFFE1;
        rom[217][62] = 16'h000C;
        rom[217][63] = 16'h0031;
        rom[217][64] = 16'hFFE1;
        rom[217][65] = 16'hFFF8;
        rom[217][66] = 16'h0013;
        rom[217][67] = 16'hFFF8;
        rom[217][68] = 16'h0005;
        rom[217][69] = 16'hFFF1;
        rom[217][70] = 16'hFFE9;
        rom[217][71] = 16'h0029;
        rom[217][72] = 16'hFFD5;
        rom[217][73] = 16'hFFF5;
        rom[217][74] = 16'h0005;
        rom[217][75] = 16'hFFAB;
        rom[217][76] = 16'hFFFD;
        rom[217][77] = 16'hFFFE;
        rom[217][78] = 16'h0014;
        rom[217][79] = 16'hFFDA;
        rom[217][80] = 16'hFFEF;
        rom[217][81] = 16'h000C;
        rom[217][82] = 16'hFFF6;
        rom[217][83] = 16'hFFCE;
        rom[217][84] = 16'hFFFC;
        rom[217][85] = 16'h0041;
        rom[217][86] = 16'hFFE7;
        rom[217][87] = 16'hFFFF;
        rom[217][88] = 16'hFFF9;
        rom[217][89] = 16'h001C;
        rom[217][90] = 16'hFFD2;
        rom[217][91] = 16'hFFF9;
        rom[217][92] = 16'hFFD5;
        rom[217][93] = 16'h0038;
        rom[217][94] = 16'hFFDC;
        rom[217][95] = 16'h000D;
        rom[217][96] = 16'h002A;
        rom[217][97] = 16'h001A;
        rom[217][98] = 16'h000C;
        rom[217][99] = 16'h0029;
        rom[217][100] = 16'hFFF6;
        rom[217][101] = 16'h0005;
        rom[217][102] = 16'h0011;
        rom[217][103] = 16'h0002;
        rom[217][104] = 16'h0004;
        rom[217][105] = 16'h0011;
        rom[217][106] = 16'hFFE6;
        rom[217][107] = 16'h0013;
        rom[217][108] = 16'hFFBC;
        rom[217][109] = 16'h002E;
        rom[217][110] = 16'hFFE1;
        rom[217][111] = 16'h0006;
        rom[217][112] = 16'hFFE2;
        rom[217][113] = 16'hFFD8;
        rom[217][114] = 16'hFFFA;
        rom[217][115] = 16'h0007;
        rom[217][116] = 16'hFFB2;
        rom[217][117] = 16'h0013;
        rom[217][118] = 16'hFFFB;
        rom[217][119] = 16'h0009;
        rom[217][120] = 16'h000E;
        rom[217][121] = 16'hFFE4;
        rom[217][122] = 16'hFFE0;
        rom[217][123] = 16'hFFE3;
        rom[217][124] = 16'h0019;
        rom[217][125] = 16'h001C;
        rom[217][126] = 16'h000D;
        rom[217][127] = 16'h0016;
        rom[218][0] = 16'hFFCD;
        rom[218][1] = 16'h000C;
        rom[218][2] = 16'hFFF9;
        rom[218][3] = 16'hFFCC;
        rom[218][4] = 16'hFFB8;
        rom[218][5] = 16'h001B;
        rom[218][6] = 16'h0017;
        rom[218][7] = 16'h0007;
        rom[218][8] = 16'h0004;
        rom[218][9] = 16'hFFD2;
        rom[218][10] = 16'h0007;
        rom[218][11] = 16'hFFEE;
        rom[218][12] = 16'h002E;
        rom[218][13] = 16'hFFF3;
        rom[218][14] = 16'hFFC3;
        rom[218][15] = 16'hFFEA;
        rom[218][16] = 16'h001E;
        rom[218][17] = 16'h0002;
        rom[218][18] = 16'hFFE6;
        rom[218][19] = 16'h0016;
        rom[218][20] = 16'h0014;
        rom[218][21] = 16'hFFF7;
        rom[218][22] = 16'h000C;
        rom[218][23] = 16'hFFD2;
        rom[218][24] = 16'hFFE4;
        rom[218][25] = 16'h001E;
        rom[218][26] = 16'hFFBC;
        rom[218][27] = 16'hFFB6;
        rom[218][28] = 16'hFFD1;
        rom[218][29] = 16'h0012;
        rom[218][30] = 16'hFFEC;
        rom[218][31] = 16'h001F;
        rom[218][32] = 16'h0007;
        rom[218][33] = 16'h0002;
        rom[218][34] = 16'h0002;
        rom[218][35] = 16'hFFE8;
        rom[218][36] = 16'h0020;
        rom[218][37] = 16'h0007;
        rom[218][38] = 16'hFFFA;
        rom[218][39] = 16'hFFF9;
        rom[218][40] = 16'hFFF3;
        rom[218][41] = 16'h000F;
        rom[218][42] = 16'hFFEF;
        rom[218][43] = 16'h0000;
        rom[218][44] = 16'hFFFF;
        rom[218][45] = 16'hFFF9;
        rom[218][46] = 16'hFFE7;
        rom[218][47] = 16'h0023;
        rom[218][48] = 16'h0029;
        rom[218][49] = 16'h0024;
        rom[218][50] = 16'h000F;
        rom[218][51] = 16'h000A;
        rom[218][52] = 16'hFFF5;
        rom[218][53] = 16'h0011;
        rom[218][54] = 16'hFFED;
        rom[218][55] = 16'hFFF2;
        rom[218][56] = 16'hFFF5;
        rom[218][57] = 16'h000E;
        rom[218][58] = 16'hFFF1;
        rom[218][59] = 16'hFFC7;
        rom[218][60] = 16'h0002;
        rom[218][61] = 16'h0010;
        rom[218][62] = 16'hFFFF;
        rom[218][63] = 16'h0033;
        rom[218][64] = 16'hFFE7;
        rom[218][65] = 16'h0026;
        rom[218][66] = 16'h0007;
        rom[218][67] = 16'h001F;
        rom[218][68] = 16'h0008;
        rom[218][69] = 16'hFFF3;
        rom[218][70] = 16'hFFFE;
        rom[218][71] = 16'h0003;
        rom[218][72] = 16'hFFD7;
        rom[218][73] = 16'hFFFF;
        rom[218][74] = 16'h0035;
        rom[218][75] = 16'hFFF3;
        rom[218][76] = 16'hFFE1;
        rom[218][77] = 16'h0016;
        rom[218][78] = 16'hFFF9;
        rom[218][79] = 16'hFFF3;
        rom[218][80] = 16'h002A;
        rom[218][81] = 16'h000F;
        rom[218][82] = 16'h001E;
        rom[218][83] = 16'hFFEF;
        rom[218][84] = 16'h0027;
        rom[218][85] = 16'h001E;
        rom[218][86] = 16'hFFCD;
        rom[218][87] = 16'h0016;
        rom[218][88] = 16'hFFFB;
        rom[218][89] = 16'h000F;
        rom[218][90] = 16'h0039;
        rom[218][91] = 16'hFFDA;
        rom[218][92] = 16'hFFD6;
        rom[218][93] = 16'hFFEA;
        rom[218][94] = 16'hFFB1;
        rom[218][95] = 16'hFFF4;
        rom[218][96] = 16'h0028;
        rom[218][97] = 16'hFFEF;
        rom[218][98] = 16'hFFEA;
        rom[218][99] = 16'hFFF0;
        rom[218][100] = 16'hFFF6;
        rom[218][101] = 16'hFFE7;
        rom[218][102] = 16'h0000;
        rom[218][103] = 16'hFFE5;
        rom[218][104] = 16'h0012;
        rom[218][105] = 16'hFFEB;
        rom[218][106] = 16'hFFF6;
        rom[218][107] = 16'h0014;
        rom[218][108] = 16'hFFD7;
        rom[218][109] = 16'hFFF9;
        rom[218][110] = 16'h0008;
        rom[218][111] = 16'h0010;
        rom[218][112] = 16'h0003;
        rom[218][113] = 16'hFFF9;
        rom[218][114] = 16'hFFD1;
        rom[218][115] = 16'h001A;
        rom[218][116] = 16'hFFEA;
        rom[218][117] = 16'h0016;
        rom[218][118] = 16'h0027;
        rom[218][119] = 16'hFFF7;
        rom[218][120] = 16'h000C;
        rom[218][121] = 16'hFFDC;
        rom[218][122] = 16'hFFCF;
        rom[218][123] = 16'hFFFC;
        rom[218][124] = 16'hFFF3;
        rom[218][125] = 16'hFFFB;
        rom[218][126] = 16'h000C;
        rom[218][127] = 16'hFFE4;
        rom[219][0] = 16'hFFE5;
        rom[219][1] = 16'hFFC0;
        rom[219][2] = 16'h0008;
        rom[219][3] = 16'hFFFB;
        rom[219][4] = 16'h000A;
        rom[219][5] = 16'hFFD6;
        rom[219][6] = 16'hFFDE;
        rom[219][7] = 16'hFFD3;
        rom[219][8] = 16'hFFAF;
        rom[219][9] = 16'h000C;
        rom[219][10] = 16'hFFE8;
        rom[219][11] = 16'h0009;
        rom[219][12] = 16'hFFEA;
        rom[219][13] = 16'hFFED;
        rom[219][14] = 16'hFFD5;
        rom[219][15] = 16'hFFD5;
        rom[219][16] = 16'hFFE3;
        rom[219][17] = 16'hFFF9;
        rom[219][18] = 16'hFFFF;
        rom[219][19] = 16'hFFF8;
        rom[219][20] = 16'h001C;
        rom[219][21] = 16'hFFD3;
        rom[219][22] = 16'hFFFC;
        rom[219][23] = 16'hFFF6;
        rom[219][24] = 16'h0003;
        rom[219][25] = 16'h0003;
        rom[219][26] = 16'hFFFB;
        rom[219][27] = 16'h0023;
        rom[219][28] = 16'h0014;
        rom[219][29] = 16'hFFC6;
        rom[219][30] = 16'hFFE9;
        rom[219][31] = 16'hFFE1;
        rom[219][32] = 16'h0002;
        rom[219][33] = 16'hFFCD;
        rom[219][34] = 16'hFFE1;
        rom[219][35] = 16'hFFD4;
        rom[219][36] = 16'hFFFB;
        rom[219][37] = 16'hFFEF;
        rom[219][38] = 16'h0009;
        rom[219][39] = 16'hFFC5;
        rom[219][40] = 16'hFF98;
        rom[219][41] = 16'hFFCF;
        rom[219][42] = 16'hFFDA;
        rom[219][43] = 16'h0027;
        rom[219][44] = 16'hFFCF;
        rom[219][45] = 16'h001A;
        rom[219][46] = 16'h000D;
        rom[219][47] = 16'h0000;
        rom[219][48] = 16'h001E;
        rom[219][49] = 16'hFFF7;
        rom[219][50] = 16'h0010;
        rom[219][51] = 16'hFFEE;
        rom[219][52] = 16'hFFE8;
        rom[219][53] = 16'h000B;
        rom[219][54] = 16'h0026;
        rom[219][55] = 16'hFFD2;
        rom[219][56] = 16'hFFD8;
        rom[219][57] = 16'h001A;
        rom[219][58] = 16'hFFEF;
        rom[219][59] = 16'h002B;
        rom[219][60] = 16'hFFE4;
        rom[219][61] = 16'hFFD7;
        rom[219][62] = 16'hFFFC;
        rom[219][63] = 16'hFFF9;
        rom[219][64] = 16'hFFE2;
        rom[219][65] = 16'hFFF1;
        rom[219][66] = 16'hFFD9;
        rom[219][67] = 16'hFFF0;
        rom[219][68] = 16'hFFCD;
        rom[219][69] = 16'hFFFC;
        rom[219][70] = 16'hFFDF;
        rom[219][71] = 16'h0006;
        rom[219][72] = 16'h000C;
        rom[219][73] = 16'hFFE8;
        rom[219][74] = 16'hFFC4;
        rom[219][75] = 16'hFFE4;
        rom[219][76] = 16'h001A;
        rom[219][77] = 16'hFFF4;
        rom[219][78] = 16'hFFC5;
        rom[219][79] = 16'hFFE7;
        rom[219][80] = 16'h0007;
        rom[219][81] = 16'h0003;
        rom[219][82] = 16'h002F;
        rom[219][83] = 16'hFFDA;
        rom[219][84] = 16'hFFF7;
        rom[219][85] = 16'h003D;
        rom[219][86] = 16'hFFF1;
        rom[219][87] = 16'h0008;
        rom[219][88] = 16'h0008;
        rom[219][89] = 16'h000C;
        rom[219][90] = 16'h0031;
        rom[219][91] = 16'hFFEF;
        rom[219][92] = 16'hFFF7;
        rom[219][93] = 16'h0008;
        rom[219][94] = 16'hFFC3;
        rom[219][95] = 16'h0002;
        rom[219][96] = 16'hFFF9;
        rom[219][97] = 16'h0000;
        rom[219][98] = 16'hFFE0;
        rom[219][99] = 16'hFFF2;
        rom[219][100] = 16'h000A;
        rom[219][101] = 16'hFFCF;
        rom[219][102] = 16'h0016;
        rom[219][103] = 16'hFFFE;
        rom[219][104] = 16'h000C;
        rom[219][105] = 16'hFFFA;
        rom[219][106] = 16'hFFE0;
        rom[219][107] = 16'h0000;
        rom[219][108] = 16'h000C;
        rom[219][109] = 16'h002A;
        rom[219][110] = 16'hFFDC;
        rom[219][111] = 16'h000C;
        rom[219][112] = 16'h0006;
        rom[219][113] = 16'hFFFE;
        rom[219][114] = 16'hFFFE;
        rom[219][115] = 16'hFFCB;
        rom[219][116] = 16'hFFE9;
        rom[219][117] = 16'hFFD6;
        rom[219][118] = 16'h0019;
        rom[219][119] = 16'h000E;
        rom[219][120] = 16'hFFFF;
        rom[219][121] = 16'hFFF9;
        rom[219][122] = 16'h0002;
        rom[219][123] = 16'hFFF6;
        rom[219][124] = 16'h001E;
        rom[219][125] = 16'h0002;
        rom[219][126] = 16'h0016;
        rom[219][127] = 16'hFFF0;
        rom[220][0] = 16'hFFE1;
        rom[220][1] = 16'h002A;
        rom[220][2] = 16'hFFE4;
        rom[220][3] = 16'hFFD2;
        rom[220][4] = 16'h000D;
        rom[220][5] = 16'h0015;
        rom[220][6] = 16'h000A;
        rom[220][7] = 16'hFFFD;
        rom[220][8] = 16'h0011;
        rom[220][9] = 16'h0002;
        rom[220][10] = 16'hFFDD;
        rom[220][11] = 16'hFFEC;
        rom[220][12] = 16'hFFEF;
        rom[220][13] = 16'hFFEA;
        rom[220][14] = 16'hFFF5;
        rom[220][15] = 16'hFFF4;
        rom[220][16] = 16'h0012;
        rom[220][17] = 16'hFFE1;
        rom[220][18] = 16'hFFE2;
        rom[220][19] = 16'h0011;
        rom[220][20] = 16'h0036;
        rom[220][21] = 16'h001D;
        rom[220][22] = 16'hFFD1;
        rom[220][23] = 16'hFFD7;
        rom[220][24] = 16'hFFED;
        rom[220][25] = 16'h001B;
        rom[220][26] = 16'h004C;
        rom[220][27] = 16'hFFD9;
        rom[220][28] = 16'h0001;
        rom[220][29] = 16'hFFF8;
        rom[220][30] = 16'hFFFF;
        rom[220][31] = 16'h0018;
        rom[220][32] = 16'hFFBF;
        rom[220][33] = 16'h001A;
        rom[220][34] = 16'hFFDD;
        rom[220][35] = 16'h000D;
        rom[220][36] = 16'h001B;
        rom[220][37] = 16'h0051;
        rom[220][38] = 16'hFFD4;
        rom[220][39] = 16'hFFF5;
        rom[220][40] = 16'hFFF4;
        rom[220][41] = 16'h001F;
        rom[220][42] = 16'hFFEE;
        rom[220][43] = 16'hFFE8;
        rom[220][44] = 16'hFFF2;
        rom[220][45] = 16'h002A;
        rom[220][46] = 16'h0010;
        rom[220][47] = 16'hFFEE;
        rom[220][48] = 16'hFFE8;
        rom[220][49] = 16'hFFFF;
        rom[220][50] = 16'hFFEC;
        rom[220][51] = 16'h0008;
        rom[220][52] = 16'hFFF4;
        rom[220][53] = 16'hFFDC;
        rom[220][54] = 16'h0007;
        rom[220][55] = 16'h0005;
        rom[220][56] = 16'hFFE0;
        rom[220][57] = 16'hFFE5;
        rom[220][58] = 16'h0008;
        rom[220][59] = 16'hFFCD;
        rom[220][60] = 16'h0007;
        rom[220][61] = 16'hFFCA;
        rom[220][62] = 16'h003B;
        rom[220][63] = 16'h0005;
        rom[220][64] = 16'hFFE2;
        rom[220][65] = 16'h0029;
        rom[220][66] = 16'h0012;
        rom[220][67] = 16'hFFFA;
        rom[220][68] = 16'h002A;
        rom[220][69] = 16'h001D;
        rom[220][70] = 16'h0010;
        rom[220][71] = 16'h0001;
        rom[220][72] = 16'h0000;
        rom[220][73] = 16'hFFE8;
        rom[220][74] = 16'h001A;
        rom[220][75] = 16'hFFE6;
        rom[220][76] = 16'hFFC8;
        rom[220][77] = 16'hFFD7;
        rom[220][78] = 16'h0007;
        rom[220][79] = 16'h0015;
        rom[220][80] = 16'h0028;
        rom[220][81] = 16'h001B;
        rom[220][82] = 16'h000A;
        rom[220][83] = 16'h0011;
        rom[220][84] = 16'hFFF7;
        rom[220][85] = 16'hFFF5;
        rom[220][86] = 16'hFFCA;
        rom[220][87] = 16'hFFFE;
        rom[220][88] = 16'h0033;
        rom[220][89] = 16'h000F;
        rom[220][90] = 16'h000A;
        rom[220][91] = 16'h0012;
        rom[220][92] = 16'h001E;
        rom[220][93] = 16'hFFDB;
        rom[220][94] = 16'hFFDE;
        rom[220][95] = 16'hFFFE;
        rom[220][96] = 16'h0018;
        rom[220][97] = 16'h0015;
        rom[220][98] = 16'hFFF7;
        rom[220][99] = 16'h0006;
        rom[220][100] = 16'hFFFE;
        rom[220][101] = 16'hFFE8;
        rom[220][102] = 16'h000A;
        rom[220][103] = 16'hFFD1;
        rom[220][104] = 16'h001A;
        rom[220][105] = 16'hFFFE;
        rom[220][106] = 16'hFFEA;
        rom[220][107] = 16'hFFDF;
        rom[220][108] = 16'hFFE8;
        rom[220][109] = 16'hFFED;
        rom[220][110] = 16'h0017;
        rom[220][111] = 16'h0005;
        rom[220][112] = 16'h000C;
        rom[220][113] = 16'hFFF7;
        rom[220][114] = 16'h0000;
        rom[220][115] = 16'h0024;
        rom[220][116] = 16'hFFF1;
        rom[220][117] = 16'h0017;
        rom[220][118] = 16'h000B;
        rom[220][119] = 16'h000D;
        rom[220][120] = 16'hFFCC;
        rom[220][121] = 16'hFFE0;
        rom[220][122] = 16'hFFC8;
        rom[220][123] = 16'hFFEA;
        rom[220][124] = 16'h0020;
        rom[220][125] = 16'hFFE1;
        rom[220][126] = 16'h0014;
        rom[220][127] = 16'h000A;
        rom[221][0] = 16'h0025;
        rom[221][1] = 16'hFFEA;
        rom[221][2] = 16'h002A;
        rom[221][3] = 16'h002E;
        rom[221][4] = 16'h001B;
        rom[221][5] = 16'hFFE3;
        rom[221][6] = 16'h002C;
        rom[221][7] = 16'hFFDE;
        rom[221][8] = 16'hFFF7;
        rom[221][9] = 16'h002F;
        rom[221][10] = 16'hFFA6;
        rom[221][11] = 16'h0009;
        rom[221][12] = 16'hFFE6;
        rom[221][13] = 16'hFFCD;
        rom[221][14] = 16'h0004;
        rom[221][15] = 16'h0017;
        rom[221][16] = 16'h000C;
        rom[221][17] = 16'hFFA4;
        rom[221][18] = 16'hFFF6;
        rom[221][19] = 16'hFFE1;
        rom[221][20] = 16'h0016;
        rom[221][21] = 16'h0016;
        rom[221][22] = 16'h001A;
        rom[221][23] = 16'hFFDA;
        rom[221][24] = 16'h0006;
        rom[221][25] = 16'h0023;
        rom[221][26] = 16'hFFF8;
        rom[221][27] = 16'hFFFF;
        rom[221][28] = 16'h0025;
        rom[221][29] = 16'h0022;
        rom[221][30] = 16'hFFFE;
        rom[221][31] = 16'h001C;
        rom[221][32] = 16'hFFFE;
        rom[221][33] = 16'hFFDD;
        rom[221][34] = 16'h0046;
        rom[221][35] = 16'h000F;
        rom[221][36] = 16'h0022;
        rom[221][37] = 16'h0004;
        rom[221][38] = 16'hFFE6;
        rom[221][39] = 16'hFFFF;
        rom[221][40] = 16'h000C;
        rom[221][41] = 16'h000C;
        rom[221][42] = 16'h0017;
        rom[221][43] = 16'hFFE4;
        rom[221][44] = 16'h0019;
        rom[221][45] = 16'hFFFF;
        rom[221][46] = 16'hFFE6;
        rom[221][47] = 16'hFFDC;
        rom[221][48] = 16'hFFF2;
        rom[221][49] = 16'hFFEA;
        rom[221][50] = 16'hFFE8;
        rom[221][51] = 16'hFFDB;
        rom[221][52] = 16'hFFFF;
        rom[221][53] = 16'hFFF4;
        rom[221][54] = 16'h0002;
        rom[221][55] = 16'hFFEE;
        rom[221][56] = 16'h0010;
        rom[221][57] = 16'h000C;
        rom[221][58] = 16'hFFB6;
        rom[221][59] = 16'h0001;
        rom[221][60] = 16'h0023;
        rom[221][61] = 16'hFFD5;
        rom[221][62] = 16'hFFF1;
        rom[221][63] = 16'h000A;
        rom[221][64] = 16'h0028;
        rom[221][65] = 16'hFFE7;
        rom[221][66] = 16'hFFF9;
        rom[221][67] = 16'hFFF5;
        rom[221][68] = 16'hFFF0;
        rom[221][69] = 16'hFFFC;
        rom[221][70] = 16'hFFFF;
        rom[221][71] = 16'h0014;
        rom[221][72] = 16'hFFF2;
        rom[221][73] = 16'hFFDB;
        rom[221][74] = 16'hFFD2;
        rom[221][75] = 16'hFFFE;
        rom[221][76] = 16'h002A;
        rom[221][77] = 16'hFFBC;
        rom[221][78] = 16'hFFFE;
        rom[221][79] = 16'hFFF4;
        rom[221][80] = 16'h0033;
        rom[221][81] = 16'hFFF7;
        rom[221][82] = 16'hFFE9;
        rom[221][83] = 16'hFFD9;
        rom[221][84] = 16'h0010;
        rom[221][85] = 16'h0013;
        rom[221][86] = 16'h0002;
        rom[221][87] = 16'h0000;
        rom[221][88] = 16'h0016;
        rom[221][89] = 16'hFFBF;
        rom[221][90] = 16'hFFF3;
        rom[221][91] = 16'h0033;
        rom[221][92] = 16'hFFFE;
        rom[221][93] = 16'h001C;
        rom[221][94] = 16'h0002;
        rom[221][95] = 16'h000E;
        rom[221][96] = 16'hFFEF;
        rom[221][97] = 16'h0003;
        rom[221][98] = 16'h0004;
        rom[221][99] = 16'hFFD8;
        rom[221][100] = 16'h000A;
        rom[221][101] = 16'h002C;
        rom[221][102] = 16'hFFE4;
        rom[221][103] = 16'h0016;
        rom[221][104] = 16'hFFF8;
        rom[221][105] = 16'h0003;
        rom[221][106] = 16'h0016;
        rom[221][107] = 16'hFFDC;
        rom[221][108] = 16'hFFD0;
        rom[221][109] = 16'h0027;
        rom[221][110] = 16'h0012;
        rom[221][111] = 16'hFFEF;
        rom[221][112] = 16'hFFF6;
        rom[221][113] = 16'h000C;
        rom[221][114] = 16'hFFE8;
        rom[221][115] = 16'h0031;
        rom[221][116] = 16'h001B;
        rom[221][117] = 16'hFFFE;
        rom[221][118] = 16'hFFFA;
        rom[221][119] = 16'hFFDD;
        rom[221][120] = 16'hFFF7;
        rom[221][121] = 16'h000A;
        rom[221][122] = 16'h0016;
        rom[221][123] = 16'hFFF8;
        rom[221][124] = 16'hFFFD;
        rom[221][125] = 16'hFFED;
        rom[221][126] = 16'h0035;
        rom[221][127] = 16'h0002;
        rom[222][0] = 16'hFFFA;
        rom[222][1] = 16'hFFFB;
        rom[222][2] = 16'h0024;
        rom[222][3] = 16'h000F;
        rom[222][4] = 16'hFFC0;
        rom[222][5] = 16'hFFF4;
        rom[222][6] = 16'hFFD5;
        rom[222][7] = 16'h0012;
        rom[222][8] = 16'h0019;
        rom[222][9] = 16'hFFFD;
        rom[222][10] = 16'hFFFE;
        rom[222][11] = 16'hFFE0;
        rom[222][12] = 16'hFFF5;
        rom[222][13] = 16'h0007;
        rom[222][14] = 16'hFFDE;
        rom[222][15] = 16'h0011;
        rom[222][16] = 16'h0006;
        rom[222][17] = 16'h0006;
        rom[222][18] = 16'hFFF3;
        rom[222][19] = 16'hFFDE;
        rom[222][20] = 16'hFFDC;
        rom[222][21] = 16'h0021;
        rom[222][22] = 16'h001E;
        rom[222][23] = 16'hFFE4;
        rom[222][24] = 16'hFFF2;
        rom[222][25] = 16'hFFD0;
        rom[222][26] = 16'hFFE1;
        rom[222][27] = 16'hFFBB;
        rom[222][28] = 16'h0012;
        rom[222][29] = 16'hFFE2;
        rom[222][30] = 16'hFFDB;
        rom[222][31] = 16'h001A;
        rom[222][32] = 16'h001B;
        rom[222][33] = 16'h0029;
        rom[222][34] = 16'h0029;
        rom[222][35] = 16'h000B;
        rom[222][36] = 16'h0014;
        rom[222][37] = 16'hFFF8;
        rom[222][38] = 16'h0013;
        rom[222][39] = 16'h0004;
        rom[222][40] = 16'hFFEA;
        rom[222][41] = 16'hFFFF;
        rom[222][42] = 16'hFFDB;
        rom[222][43] = 16'h0023;
        rom[222][44] = 16'hFFF0;
        rom[222][45] = 16'h000C;
        rom[222][46] = 16'hFFF8;
        rom[222][47] = 16'hFFD8;
        rom[222][48] = 16'h000C;
        rom[222][49] = 16'h0017;
        rom[222][50] = 16'hFFF4;
        rom[222][51] = 16'hFFF9;
        rom[222][52] = 16'h0021;
        rom[222][53] = 16'hFFEC;
        rom[222][54] = 16'hFFEB;
        rom[222][55] = 16'h0000;
        rom[222][56] = 16'h000B;
        rom[222][57] = 16'hFFC4;
        rom[222][58] = 16'h0029;
        rom[222][59] = 16'hFFD6;
        rom[222][60] = 16'hFFD9;
        rom[222][61] = 16'hFFEA;
        rom[222][62] = 16'h0007;
        rom[222][63] = 16'hFFF7;
        rom[222][64] = 16'hFFDC;
        rom[222][65] = 16'h0012;
        rom[222][66] = 16'hFFE6;
        rom[222][67] = 16'hFFE6;
        rom[222][68] = 16'hFFCD;
        rom[222][69] = 16'hFFF4;
        rom[222][70] = 16'h000E;
        rom[222][71] = 16'h0038;
        rom[222][72] = 16'hFFFE;
        rom[222][73] = 16'hFFEB;
        rom[222][74] = 16'hFFEF;
        rom[222][75] = 16'hFFEB;
        rom[222][76] = 16'h0010;
        rom[222][77] = 16'hFFE0;
        rom[222][78] = 16'h000C;
        rom[222][79] = 16'hFFDC;
        rom[222][80] = 16'hFFFF;
        rom[222][81] = 16'h001F;
        rom[222][82] = 16'hFFDB;
        rom[222][83] = 16'h001C;
        rom[222][84] = 16'h0016;
        rom[222][85] = 16'h0000;
        rom[222][86] = 16'h0013;
        rom[222][87] = 16'h000A;
        rom[222][88] = 16'hFFFE;
        rom[222][89] = 16'h000C;
        rom[222][90] = 16'hFFE4;
        rom[222][91] = 16'h0027;
        rom[222][92] = 16'h000F;
        rom[222][93] = 16'h0015;
        rom[222][94] = 16'h0007;
        rom[222][95] = 16'hFFFB;
        rom[222][96] = 16'h000C;
        rom[222][97] = 16'hFFC1;
        rom[222][98] = 16'hFFEA;
        rom[222][99] = 16'h0022;
        rom[222][100] = 16'hFFDC;
        rom[222][101] = 16'h000E;
        rom[222][102] = 16'hFFE4;
        rom[222][103] = 16'hFFD9;
        rom[222][104] = 16'hFFD3;
        rom[222][105] = 16'hFFDC;
        rom[222][106] = 16'hFFDB;
        rom[222][107] = 16'h0029;
        rom[222][108] = 16'h000B;
        rom[222][109] = 16'hFFD0;
        rom[222][110] = 16'hFFDC;
        rom[222][111] = 16'h0035;
        rom[222][112] = 16'hFFDB;
        rom[222][113] = 16'hFFCF;
        rom[222][114] = 16'hFFD2;
        rom[222][115] = 16'hFFFC;
        rom[222][116] = 16'h001D;
        rom[222][117] = 16'hFFEE;
        rom[222][118] = 16'hFFE3;
        rom[222][119] = 16'h0021;
        rom[222][120] = 16'h000B;
        rom[222][121] = 16'hFFCD;
        rom[222][122] = 16'hFFF4;
        rom[222][123] = 16'h000D;
        rom[222][124] = 16'h001F;
        rom[222][125] = 16'hFFD6;
        rom[222][126] = 16'h0024;
        rom[222][127] = 16'h0036;
        rom[223][0] = 16'hFFF1;
        rom[223][1] = 16'h0006;
        rom[223][2] = 16'hFFEF;
        rom[223][3] = 16'hFFC1;
        rom[223][4] = 16'hFFDA;
        rom[223][5] = 16'h001E;
        rom[223][6] = 16'hFFFF;
        rom[223][7] = 16'hFFF4;
        rom[223][8] = 16'h0008;
        rom[223][9] = 16'hFFC2;
        rom[223][10] = 16'hFFEA;
        rom[223][11] = 16'hFFFD;
        rom[223][12] = 16'h0008;
        rom[223][13] = 16'hFFEA;
        rom[223][14] = 16'hFFEF;
        rom[223][15] = 16'hFFF8;
        rom[223][16] = 16'h0002;
        rom[223][17] = 16'hFFE8;
        rom[223][18] = 16'hFFFE;
        rom[223][19] = 16'h0004;
        rom[223][20] = 16'h003D;
        rom[223][21] = 16'hFFD8;
        rom[223][22] = 16'hFFEA;
        rom[223][23] = 16'hFFE1;
        rom[223][24] = 16'hFFEB;
        rom[223][25] = 16'h0018;
        rom[223][26] = 16'h0015;
        rom[223][27] = 16'hFFF1;
        rom[223][28] = 16'h0000;
        rom[223][29] = 16'hFFF9;
        rom[223][30] = 16'h000D;
        rom[223][31] = 16'hFFED;
        rom[223][32] = 16'h0014;
        rom[223][33] = 16'hFFD0;
        rom[223][34] = 16'hFFC0;
        rom[223][35] = 16'hFFF7;
        rom[223][36] = 16'h000C;
        rom[223][37] = 16'h001B;
        rom[223][38] = 16'hFFFE;
        rom[223][39] = 16'h0018;
        rom[223][40] = 16'hFFDC;
        rom[223][41] = 16'h000A;
        rom[223][42] = 16'h0005;
        rom[223][43] = 16'hFFF1;
        rom[223][44] = 16'h000A;
        rom[223][45] = 16'hFFF8;
        rom[223][46] = 16'h0028;
        rom[223][47] = 16'h0024;
        rom[223][48] = 16'h0031;
        rom[223][49] = 16'hFFE3;
        rom[223][50] = 16'hFFEA;
        rom[223][51] = 16'hFFF9;
        rom[223][52] = 16'hFFCB;
        rom[223][53] = 16'hFFC6;
        rom[223][54] = 16'h0018;
        rom[223][55] = 16'hFFF7;
        rom[223][56] = 16'h000C;
        rom[223][57] = 16'h001A;
        rom[223][58] = 16'hFFEF;
        rom[223][59] = 16'hFFF6;
        rom[223][60] = 16'h0006;
        rom[223][61] = 16'h0007;
        rom[223][62] = 16'h000C;
        rom[223][63] = 16'h0016;
        rom[223][64] = 16'hFFFE;
        rom[223][65] = 16'h002B;
        rom[223][66] = 16'hFFD9;
        rom[223][67] = 16'hFFD1;
        rom[223][68] = 16'h0007;
        rom[223][69] = 16'hFFC7;
        rom[223][70] = 16'hFFD1;
        rom[223][71] = 16'hFFE6;
        rom[223][72] = 16'hFFDF;
        rom[223][73] = 16'hFFDB;
        rom[223][74] = 16'hFFF6;
        rom[223][75] = 16'hFFBC;
        rom[223][76] = 16'hFFDC;
        rom[223][77] = 16'hFFFF;
        rom[223][78] = 16'h000E;
        rom[223][79] = 16'h0016;
        rom[223][80] = 16'h0002;
        rom[223][81] = 16'h003D;
        rom[223][82] = 16'h001B;
        rom[223][83] = 16'h001F;
        rom[223][84] = 16'h0012;
        rom[223][85] = 16'hFFE4;
        rom[223][86] = 16'hFFFE;
        rom[223][87] = 16'hFFD2;
        rom[223][88] = 16'hFFEF;
        rom[223][89] = 16'hFFFD;
        rom[223][90] = 16'h0016;
        rom[223][91] = 16'hFFFA;
        rom[223][92] = 16'h0006;
        rom[223][93] = 16'hFFF7;
        rom[223][94] = 16'h0016;
        rom[223][95] = 16'h0001;
        rom[223][96] = 16'h0017;
        rom[223][97] = 16'h0006;
        rom[223][98] = 16'hFFE1;
        rom[223][99] = 16'h0018;
        rom[223][100] = 16'hFFE5;
        rom[223][101] = 16'h002C;
        rom[223][102] = 16'h0013;
        rom[223][103] = 16'hFFD8;
        rom[223][104] = 16'hFFEA;
        rom[223][105] = 16'h0005;
        rom[223][106] = 16'hFFEF;
        rom[223][107] = 16'hFFF7;
        rom[223][108] = 16'h000F;
        rom[223][109] = 16'hFFF0;
        rom[223][110] = 16'h0020;
        rom[223][111] = 16'h0020;
        rom[223][112] = 16'h0037;
        rom[223][113] = 16'h0007;
        rom[223][114] = 16'hFFF7;
        rom[223][115] = 16'hFFFE;
        rom[223][116] = 16'hFFEE;
        rom[223][117] = 16'h001B;
        rom[223][118] = 16'h0012;
        rom[223][119] = 16'h0012;
        rom[223][120] = 16'hFFF7;
        rom[223][121] = 16'hFFE5;
        rom[223][122] = 16'hFFC9;
        rom[223][123] = 16'hFFFD;
        rom[223][124] = 16'h000C;
        rom[223][125] = 16'hFFF5;
        rom[223][126] = 16'hFFB9;
        rom[223][127] = 16'hFFD9;
        rom[224][0] = 16'h0018;
        rom[224][1] = 16'hFFEB;
        rom[224][2] = 16'h0012;
        rom[224][3] = 16'hFFD8;
        rom[224][4] = 16'hFFF6;
        rom[224][5] = 16'h0003;
        rom[224][6] = 16'h0016;
        rom[224][7] = 16'hFFEC;
        rom[224][8] = 16'hFFDF;
        rom[224][9] = 16'h001C;
        rom[224][10] = 16'h0016;
        rom[224][11] = 16'hFFE5;
        rom[224][12] = 16'h0007;
        rom[224][13] = 16'hFFD0;
        rom[224][14] = 16'h001E;
        rom[224][15] = 16'h0003;
        rom[224][16] = 16'hFFF9;
        rom[224][17] = 16'hFFDA;
        rom[224][18] = 16'hFFF1;
        rom[224][19] = 16'h0011;
        rom[224][20] = 16'h001A;
        rom[224][21] = 16'h0019;
        rom[224][22] = 16'hFFE1;
        rom[224][23] = 16'h000C;
        rom[224][24] = 16'h004E;
        rom[224][25] = 16'hFFF5;
        rom[224][26] = 16'h0002;
        rom[224][27] = 16'hFFED;
        rom[224][28] = 16'h0028;
        rom[224][29] = 16'h0011;
        rom[224][30] = 16'hFFF0;
        rom[224][31] = 16'hFFD2;
        rom[224][32] = 16'hFFE1;
        rom[224][33] = 16'hFFE3;
        rom[224][34] = 16'h0008;
        rom[224][35] = 16'hFFEB;
        rom[224][36] = 16'h000E;
        rom[224][37] = 16'h0026;
        rom[224][38] = 16'h0020;
        rom[224][39] = 16'h000D;
        rom[224][40] = 16'hFFE5;
        rom[224][41] = 16'hFFFB;
        rom[224][42] = 16'hFFDA;
        rom[224][43] = 16'hFFD1;
        rom[224][44] = 16'h0002;
        rom[224][45] = 16'hFFE2;
        rom[224][46] = 16'h0002;
        rom[224][47] = 16'hFFEC;
        rom[224][48] = 16'h0022;
        rom[224][49] = 16'h0020;
        rom[224][50] = 16'h001D;
        rom[224][51] = 16'h0000;
        rom[224][52] = 16'hFFFC;
        rom[224][53] = 16'hFFFE;
        rom[224][54] = 16'hFFD8;
        rom[224][55] = 16'hFFE7;
        rom[224][56] = 16'h0009;
        rom[224][57] = 16'h001F;
        rom[224][58] = 16'h0004;
        rom[224][59] = 16'hFFF4;
        rom[224][60] = 16'hFFBD;
        rom[224][61] = 16'h000C;
        rom[224][62] = 16'h0025;
        rom[224][63] = 16'hFFFE;
        rom[224][64] = 16'h0012;
        rom[224][65] = 16'hFFF8;
        rom[224][66] = 16'hFFFE;
        rom[224][67] = 16'hFFDE;
        rom[224][68] = 16'h0031;
        rom[224][69] = 16'hFFEF;
        rom[224][70] = 16'hFFEE;
        rom[224][71] = 16'hFFF9;
        rom[224][72] = 16'h0002;
        rom[224][73] = 16'h0018;
        rom[224][74] = 16'hFFE7;
        rom[224][75] = 16'h0041;
        rom[224][76] = 16'h0021;
        rom[224][77] = 16'hFFD7;
        rom[224][78] = 16'h0011;
        rom[224][79] = 16'h001B;
        rom[224][80] = 16'hFFEA;
        rom[224][81] = 16'hFFD2;
        rom[224][82] = 16'hFFFE;
        rom[224][83] = 16'hFFDA;
        rom[224][84] = 16'h000C;
        rom[224][85] = 16'h000C;
        rom[224][86] = 16'h0016;
        rom[224][87] = 16'h0004;
        rom[224][88] = 16'hFFFE;
        rom[224][89] = 16'hFFEF;
        rom[224][90] = 16'h0007;
        rom[224][91] = 16'hFFF5;
        rom[224][92] = 16'h0016;
        rom[224][93] = 16'hFFFC;
        rom[224][94] = 16'hFFEC;
        rom[224][95] = 16'hFFF7;
        rom[224][96] = 16'h0040;
        rom[224][97] = 16'h0011;
        rom[224][98] = 16'h0014;
        rom[224][99] = 16'hFFD3;
        rom[224][100] = 16'h0011;
        rom[224][101] = 16'h0028;
        rom[224][102] = 16'h0005;
        rom[224][103] = 16'h0007;
        rom[224][104] = 16'h0007;
        rom[224][105] = 16'hFFB3;
        rom[224][106] = 16'hFFEE;
        rom[224][107] = 16'h0003;
        rom[224][108] = 16'h0005;
        rom[224][109] = 16'hFFFF;
        rom[224][110] = 16'h0016;
        rom[224][111] = 16'h001B;
        rom[224][112] = 16'h0025;
        rom[224][113] = 16'hFFF9;
        rom[224][114] = 16'h0011;
        rom[224][115] = 16'h0019;
        rom[224][116] = 16'h001C;
        rom[224][117] = 16'h0021;
        rom[224][118] = 16'hFFCC;
        rom[224][119] = 16'h0004;
        rom[224][120] = 16'h0002;
        rom[224][121] = 16'h0016;
        rom[224][122] = 16'h0004;
        rom[224][123] = 16'hFFF5;
        rom[224][124] = 16'hFFF7;
        rom[224][125] = 16'h0012;
        rom[224][126] = 16'hFFE1;
        rom[224][127] = 16'h0011;
        rom[225][0] = 16'hFFBE;
        rom[225][1] = 16'h0009;
        rom[225][2] = 16'hFFE3;
        rom[225][3] = 16'h0002;
        rom[225][4] = 16'h0009;
        rom[225][5] = 16'h0011;
        rom[225][6] = 16'h0011;
        rom[225][7] = 16'h000A;
        rom[225][8] = 16'hFFD8;
        rom[225][9] = 16'h0023;
        rom[225][10] = 16'hFFF9;
        rom[225][11] = 16'h0001;
        rom[225][12] = 16'hFFE6;
        rom[225][13] = 16'hFFF9;
        rom[225][14] = 16'hFFEA;
        rom[225][15] = 16'h0005;
        rom[225][16] = 16'h0011;
        rom[225][17] = 16'h0011;
        rom[225][18] = 16'hFFEA;
        rom[225][19] = 16'h003B;
        rom[225][20] = 16'h001B;
        rom[225][21] = 16'hFFE9;
        rom[225][22] = 16'h001F;
        rom[225][23] = 16'hFFCB;
        rom[225][24] = 16'hFFEF;
        rom[225][25] = 16'hFFD9;
        rom[225][26] = 16'hFFF8;
        rom[225][27] = 16'h0011;
        rom[225][28] = 16'h000C;
        rom[225][29] = 16'h0029;
        rom[225][30] = 16'h0035;
        rom[225][31] = 16'h0016;
        rom[225][32] = 16'h0016;
        rom[225][33] = 16'hFFD7;
        rom[225][34] = 16'h0002;
        rom[225][35] = 16'hFFF3;
        rom[225][36] = 16'h0031;
        rom[225][37] = 16'hFFD6;
        rom[225][38] = 16'h0029;
        rom[225][39] = 16'h0005;
        rom[225][40] = 16'h0012;
        rom[225][41] = 16'hFFFC;
        rom[225][42] = 16'hFFD2;
        rom[225][43] = 16'hFFEB;
        rom[225][44] = 16'hFFFD;
        rom[225][45] = 16'hFFDC;
        rom[225][46] = 16'h001F;
        rom[225][47] = 16'h0008;
        rom[225][48] = 16'h000D;
        rom[225][49] = 16'hFFCE;
        rom[225][50] = 16'h0004;
        rom[225][51] = 16'h0011;
        rom[225][52] = 16'hFFD4;
        rom[225][53] = 16'h001B;
        rom[225][54] = 16'h0017;
        rom[225][55] = 16'hFFC9;
        rom[225][56] = 16'h000E;
        rom[225][57] = 16'hFFC7;
        rom[225][58] = 16'h0001;
        rom[225][59] = 16'h0013;
        rom[225][60] = 16'h0028;
        rom[225][61] = 16'hFFF5;
        rom[225][62] = 16'hFFE5;
        rom[225][63] = 16'h0027;
        rom[225][64] = 16'h0011;
        rom[225][65] = 16'h0011;
        rom[225][66] = 16'hFFE6;
        rom[225][67] = 16'hFFFE;
        rom[225][68] = 16'hFFE0;
        rom[225][69] = 16'hFFE4;
        rom[225][70] = 16'hFFE7;
        rom[225][71] = 16'hFFF4;
        rom[225][72] = 16'h000C;
        rom[225][73] = 16'h001C;
        rom[225][74] = 16'hFFDD;
        rom[225][75] = 16'hFFC9;
        rom[225][76] = 16'hFFF5;
        rom[225][77] = 16'h001F;
        rom[225][78] = 16'h0012;
        rom[225][79] = 16'h001D;
        rom[225][80] = 16'h0006;
        rom[225][81] = 16'hFFF4;
        rom[225][82] = 16'h0012;
        rom[225][83] = 16'hFFD7;
        rom[225][84] = 16'h000C;
        rom[225][85] = 16'h0037;
        rom[225][86] = 16'h0002;
        rom[225][87] = 16'h002A;
        rom[225][88] = 16'hFFE1;
        rom[225][89] = 16'h0013;
        rom[225][90] = 16'h000D;
        rom[225][91] = 16'h000E;
        rom[225][92] = 16'hFFEF;
        rom[225][93] = 16'hFFE3;
        rom[225][94] = 16'h001F;
        rom[225][95] = 16'hFFF5;
        rom[225][96] = 16'h002C;
        rom[225][97] = 16'hFFEA;
        rom[225][98] = 16'hFFE7;
        rom[225][99] = 16'hFFEF;
        rom[225][100] = 16'hFFD7;
        rom[225][101] = 16'h0007;
        rom[225][102] = 16'hFFFA;
        rom[225][103] = 16'hFFEB;
        rom[225][104] = 16'h0029;
        rom[225][105] = 16'h0004;
        rom[225][106] = 16'h0024;
        rom[225][107] = 16'hFFA6;
        rom[225][108] = 16'hFFB0;
        rom[225][109] = 16'hFFFC;
        rom[225][110] = 16'h0052;
        rom[225][111] = 16'hFFD9;
        rom[225][112] = 16'hFFCF;
        rom[225][113] = 16'hFFF9;
        rom[225][114] = 16'hFFED;
        rom[225][115] = 16'hFFFB;
        rom[225][116] = 16'hFFED;
        rom[225][117] = 16'hFFD1;
        rom[225][118] = 16'h0001;
        rom[225][119] = 16'hFFEF;
        rom[225][120] = 16'hFFF4;
        rom[225][121] = 16'h0020;
        rom[225][122] = 16'h0018;
        rom[225][123] = 16'hFFF4;
        rom[225][124] = 16'h0024;
        rom[225][125] = 16'h001B;
        rom[225][126] = 16'hFFC7;
        rom[225][127] = 16'hFFC8;
        rom[226][0] = 16'h0010;
        rom[226][1] = 16'hFFD5;
        rom[226][2] = 16'hFFFE;
        rom[226][3] = 16'hFFE0;
        rom[226][4] = 16'h0014;
        rom[226][5] = 16'h000E;
        rom[226][6] = 16'hFFC1;
        rom[226][7] = 16'hFFF4;
        rom[226][8] = 16'hFFDF;
        rom[226][9] = 16'hFFCF;
        rom[226][10] = 16'hFFE8;
        rom[226][11] = 16'hFFEF;
        rom[226][12] = 16'h000F;
        rom[226][13] = 16'h0018;
        rom[226][14] = 16'hFFF6;
        rom[226][15] = 16'hFFFB;
        rom[226][16] = 16'hFFD7;
        rom[226][17] = 16'hFFF3;
        rom[226][18] = 16'hFFB6;
        rom[226][19] = 16'hFFF6;
        rom[226][20] = 16'hFFB3;
        rom[226][21] = 16'hFFEF;
        rom[226][22] = 16'h000D;
        rom[226][23] = 16'hFFC1;
        rom[226][24] = 16'hFFF4;
        rom[226][25] = 16'hFFE5;
        rom[226][26] = 16'hFFD0;
        rom[226][27] = 16'hFFE9;
        rom[226][28] = 16'hFFEA;
        rom[226][29] = 16'hFFE1;
        rom[226][30] = 16'h0011;
        rom[226][31] = 16'h0016;
        rom[226][32] = 16'hFFF4;
        rom[226][33] = 16'h000F;
        rom[226][34] = 16'h0000;
        rom[226][35] = 16'h0012;
        rom[226][36] = 16'hFFE3;
        rom[226][37] = 16'hFFC8;
        rom[226][38] = 16'hFFB0;
        rom[226][39] = 16'h000D;
        rom[226][40] = 16'h0014;
        rom[226][41] = 16'hFFB6;
        rom[226][42] = 16'h000F;
        rom[226][43] = 16'hFFEF;
        rom[226][44] = 16'h0039;
        rom[226][45] = 16'h0015;
        rom[226][46] = 16'hFFAE;
        rom[226][47] = 16'h001A;
        rom[226][48] = 16'h001C;
        rom[226][49] = 16'h000D;
        rom[226][50] = 16'h0010;
        rom[226][51] = 16'h0006;
        rom[226][52] = 16'h0012;
        rom[226][53] = 16'hFFF4;
        rom[226][54] = 16'hFFE4;
        rom[226][55] = 16'hFFEA;
        rom[226][56] = 16'h0026;
        rom[226][57] = 16'h000E;
        rom[226][58] = 16'hFFFC;
        rom[226][59] = 16'hFFD7;
        rom[226][60] = 16'h0006;
        rom[226][61] = 16'h000A;
        rom[226][62] = 16'hFFDE;
        rom[226][63] = 16'h000B;
        rom[226][64] = 16'hFFC3;
        rom[226][65] = 16'hFFB0;
        rom[226][66] = 16'h0007;
        rom[226][67] = 16'hFFFD;
        rom[226][68] = 16'hFFF4;
        rom[226][69] = 16'h0005;
        rom[226][70] = 16'hFFF7;
        rom[226][71] = 16'hFFEC;
        rom[226][72] = 16'h0010;
        rom[226][73] = 16'hFFED;
        rom[226][74] = 16'hFFD8;
        rom[226][75] = 16'hFFD6;
        rom[226][76] = 16'hFFD2;
        rom[226][77] = 16'h0004;
        rom[226][78] = 16'hFFFE;
        rom[226][79] = 16'h0010;
        rom[226][80] = 16'hFFBB;
        rom[226][81] = 16'hFFFE;
        rom[226][82] = 16'hFFE3;
        rom[226][83] = 16'h0008;
        rom[226][84] = 16'h0006;
        rom[226][85] = 16'h001B;
        rom[226][86] = 16'hFFD6;
        rom[226][87] = 16'h0007;
        rom[226][88] = 16'hFFC9;
        rom[226][89] = 16'h0019;
        rom[226][90] = 16'hFFCF;
        rom[226][91] = 16'hFFC2;
        rom[226][92] = 16'hFFDC;
        rom[226][93] = 16'h0018;
        rom[226][94] = 16'hFFF4;
        rom[226][95] = 16'h0033;
        rom[226][96] = 16'h0016;
        rom[226][97] = 16'hFFEA;
        rom[226][98] = 16'hFFFB;
        rom[226][99] = 16'hFFE0;
        rom[226][100] = 16'hFFFB;
        rom[226][101] = 16'hFFE7;
        rom[226][102] = 16'hFFF2;
        rom[226][103] = 16'h0019;
        rom[226][104] = 16'h001B;
        rom[226][105] = 16'hFFFD;
        rom[226][106] = 16'hFFDB;
        rom[226][107] = 16'h0011;
        rom[226][108] = 16'hFFE2;
        rom[226][109] = 16'hFFFE;
        rom[226][110] = 16'hFFFE;
        rom[226][111] = 16'hFFE3;
        rom[226][112] = 16'h0011;
        rom[226][113] = 16'hFFFC;
        rom[226][114] = 16'h0005;
        rom[226][115] = 16'hFFE8;
        rom[226][116] = 16'hFFB3;
        rom[226][117] = 16'hFFA9;
        rom[226][118] = 16'hFFF4;
        rom[226][119] = 16'h000F;
        rom[226][120] = 16'h0009;
        rom[226][121] = 16'hFFC8;
        rom[226][122] = 16'hFFE8;
        rom[226][123] = 16'hFFD4;
        rom[226][124] = 16'hFFFA;
        rom[226][125] = 16'h0016;
        rom[226][126] = 16'h000F;
        rom[226][127] = 16'h000F;
        rom[227][0] = 16'hFFDE;
        rom[227][1] = 16'h0003;
        rom[227][2] = 16'h0009;
        rom[227][3] = 16'hFFF8;
        rom[227][4] = 16'h000A;
        rom[227][5] = 16'hFFFF;
        rom[227][6] = 16'h002C;
        rom[227][7] = 16'hFFD0;
        rom[227][8] = 16'h002A;
        rom[227][9] = 16'h0021;
        rom[227][10] = 16'hFFFE;
        rom[227][11] = 16'h001E;
        rom[227][12] = 16'hFFF4;
        rom[227][13] = 16'hFFF4;
        rom[227][14] = 16'hFFEA;
        rom[227][15] = 16'h0018;
        rom[227][16] = 16'h001B;
        rom[227][17] = 16'h0002;
        rom[227][18] = 16'hFFD6;
        rom[227][19] = 16'h0012;
        rom[227][20] = 16'hFFAB;
        rom[227][21] = 16'h0028;
        rom[227][22] = 16'h000C;
        rom[227][23] = 16'hFFFC;
        rom[227][24] = 16'h0027;
        rom[227][25] = 16'h0008;
        rom[227][26] = 16'h002E;
        rom[227][27] = 16'hFFC2;
        rom[227][28] = 16'hFFBA;
        rom[227][29] = 16'hFFD0;
        rom[227][30] = 16'hFFED;
        rom[227][31] = 16'hFFD1;
        rom[227][32] = 16'hFFEF;
        rom[227][33] = 16'hFFF7;
        rom[227][34] = 16'h0012;
        rom[227][35] = 16'hFFC9;
        rom[227][36] = 16'h001E;
        rom[227][37] = 16'h0005;
        rom[227][38] = 16'h0026;
        rom[227][39] = 16'h0033;
        rom[227][40] = 16'hFFF6;
        rom[227][41] = 16'h0038;
        rom[227][42] = 16'hFFE7;
        rom[227][43] = 16'hFFD4;
        rom[227][44] = 16'h003E;
        rom[227][45] = 16'hFFFB;
        rom[227][46] = 16'h0016;
        rom[227][47] = 16'hFFE5;
        rom[227][48] = 16'h0007;
        rom[227][49] = 16'hFFE1;
        rom[227][50] = 16'h0022;
        rom[227][51] = 16'hFFE5;
        rom[227][52] = 16'h001E;
        rom[227][53] = 16'h0007;
        rom[227][54] = 16'h0002;
        rom[227][55] = 16'h0006;
        rom[227][56] = 16'hFFFD;
        rom[227][57] = 16'h0019;
        rom[227][58] = 16'hFFF4;
        rom[227][59] = 16'hFFDB;
        rom[227][60] = 16'hFFF0;
        rom[227][61] = 16'hFFC3;
        rom[227][62] = 16'h0007;
        rom[227][63] = 16'h0010;
        rom[227][64] = 16'hFFAD;
        rom[227][65] = 16'h0002;
        rom[227][66] = 16'h001A;
        rom[227][67] = 16'h000D;
        rom[227][68] = 16'h001F;
        rom[227][69] = 16'h001F;
        rom[227][70] = 16'h001C;
        rom[227][71] = 16'hFFFA;
        rom[227][72] = 16'hFFE2;
        rom[227][73] = 16'h0000;
        rom[227][74] = 16'hFFE5;
        rom[227][75] = 16'h0014;
        rom[227][76] = 16'h0024;
        rom[227][77] = 16'h0002;
        rom[227][78] = 16'h0041;
        rom[227][79] = 16'hFFF7;
        rom[227][80] = 16'hFFEF;
        rom[227][81] = 16'h0011;
        rom[227][82] = 16'h0000;
        rom[227][83] = 16'hFFFA;
        rom[227][84] = 16'h001E;
        rom[227][85] = 16'h000C;
        rom[227][86] = 16'hFFBF;
        rom[227][87] = 16'hFFFE;
        rom[227][88] = 16'hFFE1;
        rom[227][89] = 16'hFFFE;
        rom[227][90] = 16'hFFC6;
        rom[227][91] = 16'h0016;
        rom[227][92] = 16'h002D;
        rom[227][93] = 16'hFFD1;
        rom[227][94] = 16'h0005;
        rom[227][95] = 16'hFFF8;
        rom[227][96] = 16'hFFE5;
        rom[227][97] = 16'hFFF0;
        rom[227][98] = 16'hFFFE;
        rom[227][99] = 16'hFFF2;
        rom[227][100] = 16'hFFEE;
        rom[227][101] = 16'hFFFF;
        rom[227][102] = 16'hFFDE;
        rom[227][103] = 16'hFFEA;
        rom[227][104] = 16'h0024;
        rom[227][105] = 16'h0013;
        rom[227][106] = 16'hFFF5;
        rom[227][107] = 16'h0033;
        rom[227][108] = 16'hFFD7;
        rom[227][109] = 16'hFFCC;
        rom[227][110] = 16'hFFDA;
        rom[227][111] = 16'h0001;
        rom[227][112] = 16'hFFE4;
        rom[227][113] = 16'h0022;
        rom[227][114] = 16'hFFF7;
        rom[227][115] = 16'hFFF1;
        rom[227][116] = 16'h0007;
        rom[227][117] = 16'hFFFF;
        rom[227][118] = 16'hFFD6;
        rom[227][119] = 16'hFFF9;
        rom[227][120] = 16'hFFEE;
        rom[227][121] = 16'hFFF4;
        rom[227][122] = 16'h0024;
        rom[227][123] = 16'h0032;
        rom[227][124] = 16'hFFF7;
        rom[227][125] = 16'h0007;
        rom[227][126] = 16'h0005;
        rom[227][127] = 16'h0002;
        rom[228][0] = 16'hFFF5;
        rom[228][1] = 16'hFFD0;
        rom[228][2] = 16'hFFF2;
        rom[228][3] = 16'h0007;
        rom[228][4] = 16'h000E;
        rom[228][5] = 16'hFFCC;
        rom[228][6] = 16'h0029;
        rom[228][7] = 16'hFFE1;
        rom[228][8] = 16'hFFFD;
        rom[228][9] = 16'hFFF2;
        rom[228][10] = 16'h0009;
        rom[228][11] = 16'h000E;
        rom[228][12] = 16'hFFFC;
        rom[228][13] = 16'h0016;
        rom[228][14] = 16'h000D;
        rom[228][15] = 16'hFFFD;
        rom[228][16] = 16'h0006;
        rom[228][17] = 16'hFFB0;
        rom[228][18] = 16'h000C;
        rom[228][19] = 16'hFFD8;
        rom[228][20] = 16'hFFE1;
        rom[228][21] = 16'h001F;
        rom[228][22] = 16'hFFF9;
        rom[228][23] = 16'hFFF1;
        rom[228][24] = 16'h001B;
        rom[228][25] = 16'hFFFE;
        rom[228][26] = 16'hFFDC;
        rom[228][27] = 16'h0038;
        rom[228][28] = 16'h0027;
        rom[228][29] = 16'hFFA7;
        rom[228][30] = 16'h0016;
        rom[228][31] = 16'hFFFD;
        rom[228][32] = 16'hFFEA;
        rom[228][33] = 16'h001B;
        rom[228][34] = 16'hFFFB;
        rom[228][35] = 16'h0000;
        rom[228][36] = 16'hFFEA;
        rom[228][37] = 16'h000C;
        rom[228][38] = 16'hFFFC;
        rom[228][39] = 16'hFFDD;
        rom[228][40] = 16'hFFC8;
        rom[228][41] = 16'hFFDA;
        rom[228][42] = 16'h001B;
        rom[228][43] = 16'h0016;
        rom[228][44] = 16'hFFF0;
        rom[228][45] = 16'hFFE1;
        rom[228][46] = 16'hFFF7;
        rom[228][47] = 16'hFFC4;
        rom[228][48] = 16'hFFB2;
        rom[228][49] = 16'hFFF3;
        rom[228][50] = 16'hFFEA;
        rom[228][51] = 16'hFFF6;
        rom[228][52] = 16'hFFF5;
        rom[228][53] = 16'hFFBA;
        rom[228][54] = 16'hFFF0;
        rom[228][55] = 16'hFFF4;
        rom[228][56] = 16'hFFE0;
        rom[228][57] = 16'hFFB0;
        rom[228][58] = 16'hFFFA;
        rom[228][59] = 16'hFFF8;
        rom[228][60] = 16'h0013;
        rom[228][61] = 16'h0004;
        rom[228][62] = 16'hFFF6;
        rom[228][63] = 16'hFFC3;
        rom[228][64] = 16'hFFF7;
        rom[228][65] = 16'h001E;
        rom[228][66] = 16'hFFF0;
        rom[228][67] = 16'hFFFD;
        rom[228][68] = 16'hFFDA;
        rom[228][69] = 16'hFFE5;
        rom[228][70] = 16'hFFEE;
        rom[228][71] = 16'hFFFC;
        rom[228][72] = 16'h002F;
        rom[228][73] = 16'hFFF7;
        rom[228][74] = 16'hFFC9;
        rom[228][75] = 16'h0009;
        rom[228][76] = 16'hFFF7;
        rom[228][77] = 16'h001B;
        rom[228][78] = 16'hFFC2;
        rom[228][79] = 16'h0018;
        rom[228][80] = 16'hFFE9;
        rom[228][81] = 16'hFFEE;
        rom[228][82] = 16'hFFB1;
        rom[228][83] = 16'hFFFB;
        rom[228][84] = 16'hFFFC;
        rom[228][85] = 16'h0015;
        rom[228][86] = 16'hFFD7;
        rom[228][87] = 16'h0011;
        rom[228][88] = 16'hFFE0;
        rom[228][89] = 16'hFFC9;
        rom[228][90] = 16'hFFEF;
        rom[228][91] = 16'h0038;
        rom[228][92] = 16'h0031;
        rom[228][93] = 16'h0005;
        rom[228][94] = 16'hFFDD;
        rom[228][95] = 16'h0006;
        rom[228][96] = 16'hFFBD;
        rom[228][97] = 16'h000A;
        rom[228][98] = 16'hFFFF;
        rom[228][99] = 16'h0005;
        rom[228][100] = 16'h0021;
        rom[228][101] = 16'hFFE5;
        rom[228][102] = 16'h0014;
        rom[228][103] = 16'h003C;
        rom[228][104] = 16'h0029;
        rom[228][105] = 16'hFFD5;
        rom[228][106] = 16'h0018;
        rom[228][107] = 16'h000C;
        rom[228][108] = 16'h0027;
        rom[228][109] = 16'h0001;
        rom[228][110] = 16'hFFD4;
        rom[228][111] = 16'h0016;
        rom[228][112] = 16'h001A;
        rom[228][113] = 16'h0005;
        rom[228][114] = 16'h002E;
        rom[228][115] = 16'h000B;
        rom[228][116] = 16'hFFFD;
        rom[228][117] = 16'hFFF8;
        rom[228][118] = 16'h0005;
        rom[228][119] = 16'hFFE7;
        rom[228][120] = 16'hFFFC;
        rom[228][121] = 16'h003C;
        rom[228][122] = 16'h0024;
        rom[228][123] = 16'h002C;
        rom[228][124] = 16'h0017;
        rom[228][125] = 16'h0046;
        rom[228][126] = 16'h001A;
        rom[228][127] = 16'h0012;
        rom[229][0] = 16'h0017;
        rom[229][1] = 16'h0011;
        rom[229][2] = 16'h001D;
        rom[229][3] = 16'h0006;
        rom[229][4] = 16'hFFDD;
        rom[229][5] = 16'hFFFA;
        rom[229][6] = 16'h0024;
        rom[229][7] = 16'h001E;
        rom[229][8] = 16'hFFDA;
        rom[229][9] = 16'hFFD8;
        rom[229][10] = 16'hFFF4;
        rom[229][11] = 16'hFFF4;
        rom[229][12] = 16'hFFFE;
        rom[229][13] = 16'hFFF8;
        rom[229][14] = 16'hFFED;
        rom[229][15] = 16'h000D;
        rom[229][16] = 16'h002A;
        rom[229][17] = 16'hFFE0;
        rom[229][18] = 16'hFFF9;
        rom[229][19] = 16'h0001;
        rom[229][20] = 16'hFFE9;
        rom[229][21] = 16'hFFF4;
        rom[229][22] = 16'h001C;
        rom[229][23] = 16'hFFCE;
        rom[229][24] = 16'hFFFC;
        rom[229][25] = 16'h0009;
        rom[229][26] = 16'hFFEA;
        rom[229][27] = 16'hFFFE;
        rom[229][28] = 16'h0001;
        rom[229][29] = 16'h0019;
        rom[229][30] = 16'hFFD3;
        rom[229][31] = 16'hFFD6;
        rom[229][32] = 16'hFFF8;
        rom[229][33] = 16'hFFEF;
        rom[229][34] = 16'h0014;
        rom[229][35] = 16'hFFF4;
        rom[229][36] = 16'h0021;
        rom[229][37] = 16'hFFF4;
        rom[229][38] = 16'hFFF8;
        rom[229][39] = 16'hFFFA;
        rom[229][40] = 16'hFFF9;
        rom[229][41] = 16'hFFEB;
        rom[229][42] = 16'hFFF5;
        rom[229][43] = 16'hFFE4;
        rom[229][44] = 16'h0003;
        rom[229][45] = 16'hFFFE;
        rom[229][46] = 16'h0002;
        rom[229][47] = 16'hFFD7;
        rom[229][48] = 16'hFFF4;
        rom[229][49] = 16'h0013;
        rom[229][50] = 16'h0016;
        rom[229][51] = 16'hFFE6;
        rom[229][52] = 16'h0008;
        rom[229][53] = 16'hFFDA;
        rom[229][54] = 16'h0001;
        rom[229][55] = 16'h0006;
        rom[229][56] = 16'hFFF4;
        rom[229][57] = 16'hFFD3;
        rom[229][58] = 16'h0014;
        rom[229][59] = 16'hFFD7;
        rom[229][60] = 16'h0016;
        rom[229][61] = 16'h000A;
        rom[229][62] = 16'h0004;
        rom[229][63] = 16'h0012;
        rom[229][64] = 16'h002E;
        rom[229][65] = 16'hFFEF;
        rom[229][66] = 16'hFFF8;
        rom[229][67] = 16'hFFDF;
        rom[229][68] = 16'hFFFA;
        rom[229][69] = 16'hFFF1;
        rom[229][70] = 16'h0027;
        rom[229][71] = 16'h003D;
        rom[229][72] = 16'hFFE9;
        rom[229][73] = 16'hFFEC;
        rom[229][74] = 16'hFFE1;
        rom[229][75] = 16'hFFED;
        rom[229][76] = 16'h0020;
        rom[229][77] = 16'hFFA6;
        rom[229][78] = 16'hFFEF;
        rom[229][79] = 16'hFFEA;
        rom[229][80] = 16'hFFF9;
        rom[229][81] = 16'h0029;
        rom[229][82] = 16'h0006;
        rom[229][83] = 16'hFFFC;
        rom[229][84] = 16'h0010;
        rom[229][85] = 16'hFFC3;
        rom[229][86] = 16'hFFDF;
        rom[229][87] = 16'hFFDC;
        rom[229][88] = 16'hFFE3;
        rom[229][89] = 16'hFFF2;
        rom[229][90] = 16'h0003;
        rom[229][91] = 16'h0001;
        rom[229][92] = 16'hFFED;
        rom[229][93] = 16'h002E;
        rom[229][94] = 16'hFFCE;
        rom[229][95] = 16'hFFB5;
        rom[229][96] = 16'hFFEE;
        rom[229][97] = 16'hFFF4;
        rom[229][98] = 16'h0018;
        rom[229][99] = 16'h000C;
        rom[229][100] = 16'hFFC9;
        rom[229][101] = 16'h0014;
        rom[229][102] = 16'h003E;
        rom[229][103] = 16'h000F;
        rom[229][104] = 16'hFFF4;
        rom[229][105] = 16'hFFB9;
        rom[229][106] = 16'h001F;
        rom[229][107] = 16'h0024;
        rom[229][108] = 16'hFFFD;
        rom[229][109] = 16'h003C;
        rom[229][110] = 16'h001B;
        rom[229][111] = 16'hFFF9;
        rom[229][112] = 16'hFFDC;
        rom[229][113] = 16'hFFEC;
        rom[229][114] = 16'h0033;
        rom[229][115] = 16'h001B;
        rom[229][116] = 16'h000C;
        rom[229][117] = 16'hFFC4;
        rom[229][118] = 16'hFFDA;
        rom[229][119] = 16'h001C;
        rom[229][120] = 16'hFFE1;
        rom[229][121] = 16'hFFE3;
        rom[229][122] = 16'hFFE2;
        rom[229][123] = 16'hFFEF;
        rom[229][124] = 16'h0011;
        rom[229][125] = 16'hFFB0;
        rom[229][126] = 16'hFFF5;
        rom[229][127] = 16'hFFF1;
        rom[230][0] = 16'h0005;
        rom[230][1] = 16'hFFF5;
        rom[230][2] = 16'hFFED;
        rom[230][3] = 16'hFFA4;
        rom[230][4] = 16'h001B;
        rom[230][5] = 16'h0007;
        rom[230][6] = 16'h0002;
        rom[230][7] = 16'h0007;
        rom[230][8] = 16'hFFF5;
        rom[230][9] = 16'hFFC8;
        rom[230][10] = 16'hFFF0;
        rom[230][11] = 16'hFFB1;
        rom[230][12] = 16'hFFEC;
        rom[230][13] = 16'h0033;
        rom[230][14] = 16'hFFCB;
        rom[230][15] = 16'hFFFB;
        rom[230][16] = 16'hFFEA;
        rom[230][17] = 16'h002E;
        rom[230][18] = 16'hFFDD;
        rom[230][19] = 16'hFFEF;
        rom[230][20] = 16'hFFBA;
        rom[230][21] = 16'h0006;
        rom[230][22] = 16'hFFCD;
        rom[230][23] = 16'hFFF9;
        rom[230][24] = 16'h0016;
        rom[230][25] = 16'h000B;
        rom[230][26] = 16'hFFDA;
        rom[230][27] = 16'hFFF9;
        rom[230][28] = 16'hFFCE;
        rom[230][29] = 16'hFFE7;
        rom[230][30] = 16'h0030;
        rom[230][31] = 16'h0011;
        rom[230][32] = 16'hFFE6;
        rom[230][33] = 16'h0023;
        rom[230][34] = 16'hFFE7;
        rom[230][35] = 16'hFFD4;
        rom[230][36] = 16'h0002;
        rom[230][37] = 16'hFFF6;
        rom[230][38] = 16'hFFF7;
        rom[230][39] = 16'h0008;
        rom[230][40] = 16'h000F;
        rom[230][41] = 16'h0001;
        rom[230][42] = 16'hFFC3;
        rom[230][43] = 16'hFFEF;
        rom[230][44] = 16'h003D;
        rom[230][45] = 16'hFFDA;
        rom[230][46] = 16'hFFDE;
        rom[230][47] = 16'hFFFD;
        rom[230][48] = 16'h0010;
        rom[230][49] = 16'h000D;
        rom[230][50] = 16'hFFE3;
        rom[230][51] = 16'h0039;
        rom[230][52] = 16'hFFED;
        rom[230][53] = 16'hFFF0;
        rom[230][54] = 16'hFFD1;
        rom[230][55] = 16'hFFD3;
        rom[230][56] = 16'h002E;
        rom[230][57] = 16'h001B;
        rom[230][58] = 16'h0011;
        rom[230][59] = 16'hFFB9;
        rom[230][60] = 16'h0001;
        rom[230][61] = 16'h001D;
        rom[230][62] = 16'hFFDC;
        rom[230][63] = 16'hFFFE;
        rom[230][64] = 16'h0016;
        rom[230][65] = 16'h0022;
        rom[230][66] = 16'h0019;
        rom[230][67] = 16'h0004;
        rom[230][68] = 16'h0030;
        rom[230][69] = 16'hFFF9;
        rom[230][70] = 16'hFFED;
        rom[230][71] = 16'hFFCF;
        rom[230][72] = 16'h004B;
        rom[230][73] = 16'h000D;
        rom[230][74] = 16'h001C;
        rom[230][75] = 16'h0007;
        rom[230][76] = 16'hFFE8;
        rom[230][77] = 16'h0028;
        rom[230][78] = 16'hFFD8;
        rom[230][79] = 16'hFFF5;
        rom[230][80] = 16'h0008;
        rom[230][81] = 16'hFFF7;
        rom[230][82] = 16'hFFF9;
        rom[230][83] = 16'h001B;
        rom[230][84] = 16'hFFF0;
        rom[230][85] = 16'hFFE4;
        rom[230][86] = 16'h0007;
        rom[230][87] = 16'h0010;
        rom[230][88] = 16'h0012;
        rom[230][89] = 16'h000C;
        rom[230][90] = 16'h0001;
        rom[230][91] = 16'hFFDE;
        rom[230][92] = 16'h000C;
        rom[230][93] = 16'hFFE5;
        rom[230][94] = 16'hFFF7;
        rom[230][95] = 16'hFFF3;
        rom[230][96] = 16'h0018;
        rom[230][97] = 16'h0049;
        rom[230][98] = 16'h0023;
        rom[230][99] = 16'hFFE5;
        rom[230][100] = 16'hFFD7;
        rom[230][101] = 16'hFFF9;
        rom[230][102] = 16'h0003;
        rom[230][103] = 16'hFFFF;
        rom[230][104] = 16'h003D;
        rom[230][105] = 16'h000E;
        rom[230][106] = 16'hFFE1;
        rom[230][107] = 16'hFFCB;
        rom[230][108] = 16'hFFD9;
        rom[230][109] = 16'hFFE6;
        rom[230][110] = 16'h0016;
        rom[230][111] = 16'hFFC5;
        rom[230][112] = 16'hFFBA;
        rom[230][113] = 16'hFFD2;
        rom[230][114] = 16'hFFF4;
        rom[230][115] = 16'hFFD7;
        rom[230][116] = 16'hFFED;
        rom[230][117] = 16'hFFF4;
        rom[230][118] = 16'hFFCC;
        rom[230][119] = 16'h0002;
        rom[230][120] = 16'hFFF0;
        rom[230][121] = 16'hFFD7;
        rom[230][122] = 16'hFFA7;
        rom[230][123] = 16'hFFF0;
        rom[230][124] = 16'h0003;
        rom[230][125] = 16'h001F;
        rom[230][126] = 16'hFFCB;
        rom[230][127] = 16'hFFE1;
        rom[231][0] = 16'hFFFE;
        rom[231][1] = 16'hFFCA;
        rom[231][2] = 16'hFFF1;
        rom[231][3] = 16'hFFEA;
        rom[231][4] = 16'hFFDC;
        rom[231][5] = 16'hFFD8;
        rom[231][6] = 16'h0008;
        rom[231][7] = 16'h0002;
        rom[231][8] = 16'hFFFE;
        rom[231][9] = 16'hFFFA;
        rom[231][10] = 16'h0004;
        rom[231][11] = 16'h0003;
        rom[231][12] = 16'hFFCE;
        rom[231][13] = 16'hFFC8;
        rom[231][14] = 16'h000D;
        rom[231][15] = 16'hFFD0;
        rom[231][16] = 16'h001A;
        rom[231][17] = 16'h000C;
        rom[231][18] = 16'h0017;
        rom[231][19] = 16'h0039;
        rom[231][20] = 16'hFFF7;
        rom[231][21] = 16'hFFFE;
        rom[231][22] = 16'hFFF3;
        rom[231][23] = 16'h0005;
        rom[231][24] = 16'h0003;
        rom[231][25] = 16'h0009;
        rom[231][26] = 16'hFFFD;
        rom[231][27] = 16'h0021;
        rom[231][28] = 16'h001D;
        rom[231][29] = 16'h000B;
        rom[231][30] = 16'h0002;
        rom[231][31] = 16'h0019;
        rom[231][32] = 16'h0001;
        rom[231][33] = 16'h0004;
        rom[231][34] = 16'hFFF9;
        rom[231][35] = 16'h001E;
        rom[231][36] = 16'hFFF1;
        rom[231][37] = 16'h0003;
        rom[231][38] = 16'h001A;
        rom[231][39] = 16'h002E;
        rom[231][40] = 16'hFFDC;
        rom[231][41] = 16'hFFEA;
        rom[231][42] = 16'hFFEE;
        rom[231][43] = 16'hFFE4;
        rom[231][44] = 16'hFFE4;
        rom[231][45] = 16'hFFF6;
        rom[231][46] = 16'h002D;
        rom[231][47] = 16'h0006;
        rom[231][48] = 16'hFFC2;
        rom[231][49] = 16'hFFFF;
        rom[231][50] = 16'hFFC7;
        rom[231][51] = 16'hFFE1;
        rom[231][52] = 16'hFFFC;
        rom[231][53] = 16'hFFC9;
        rom[231][54] = 16'hFFDB;
        rom[231][55] = 16'h000C;
        rom[231][56] = 16'hFFF5;
        rom[231][57] = 16'hFFF4;
        rom[231][58] = 16'hFFF7;
        rom[231][59] = 16'h001D;
        rom[231][60] = 16'hFFFD;
        rom[231][61] = 16'h002A;
        rom[231][62] = 16'h003A;
        rom[231][63] = 16'hFFF9;
        rom[231][64] = 16'hFFE5;
        rom[231][65] = 16'hFFCA;
        rom[231][66] = 16'hFFD7;
        rom[231][67] = 16'hFFEE;
        rom[231][68] = 16'hFFDA;
        rom[231][69] = 16'hFFDD;
        rom[231][70] = 16'hFFD1;
        rom[231][71] = 16'h0002;
        rom[231][72] = 16'h0010;
        rom[231][73] = 16'h0003;
        rom[231][74] = 16'hFFC5;
        rom[231][75] = 16'hFFFD;
        rom[231][76] = 16'hFFFB;
        rom[231][77] = 16'hFFDC;
        rom[231][78] = 16'hFFE5;
        rom[231][79] = 16'h0008;
        rom[231][80] = 16'h0002;
        rom[231][81] = 16'hFFEF;
        rom[231][82] = 16'hFFFE;
        rom[231][83] = 16'hFFDF;
        rom[231][84] = 16'hFFDB;
        rom[231][85] = 16'h0003;
        rom[231][86] = 16'h0039;
        rom[231][87] = 16'hFFDC;
        rom[231][88] = 16'hFFE9;
        rom[231][89] = 16'hFFEA;
        rom[231][90] = 16'h0013;
        rom[231][91] = 16'hFFE2;
        rom[231][92] = 16'hFFD7;
        rom[231][93] = 16'h001C;
        rom[231][94] = 16'hFFDE;
        rom[231][95] = 16'h0000;
        rom[231][96] = 16'hFFEF;
        rom[231][97] = 16'hFFBA;
        rom[231][98] = 16'h0000;
        rom[231][99] = 16'hFFCD;
        rom[231][100] = 16'h0018;
        rom[231][101] = 16'hFFD4;
        rom[231][102] = 16'hFFF3;
        rom[231][103] = 16'hFFDF;
        rom[231][104] = 16'hFFC5;
        rom[231][105] = 16'h0005;
        rom[231][106] = 16'hFFEE;
        rom[231][107] = 16'hFFF4;
        rom[231][108] = 16'h001B;
        rom[231][109] = 16'hFFFF;
        rom[231][110] = 16'h0029;
        rom[231][111] = 16'h0011;
        rom[231][112] = 16'hFFF9;
        rom[231][113] = 16'hFFE2;
        rom[231][114] = 16'h0002;
        rom[231][115] = 16'h0002;
        rom[231][116] = 16'h0003;
        rom[231][117] = 16'hFFF5;
        rom[231][118] = 16'hFFE4;
        rom[231][119] = 16'h0008;
        rom[231][120] = 16'hFFE0;
        rom[231][121] = 16'h001F;
        rom[231][122] = 16'hFFF9;
        rom[231][123] = 16'hFFE3;
        rom[231][124] = 16'hFFF2;
        rom[231][125] = 16'hFFD7;
        rom[231][126] = 16'h001B;
        rom[231][127] = 16'h0010;
        rom[232][0] = 16'h0024;
        rom[232][1] = 16'hFFD3;
        rom[232][2] = 16'hFFF2;
        rom[232][3] = 16'h001F;
        rom[232][4] = 16'h0008;
        rom[232][5] = 16'hFFE1;
        rom[232][6] = 16'hFFE7;
        rom[232][7] = 16'hFFD5;
        rom[232][8] = 16'hFFEF;
        rom[232][9] = 16'h000D;
        rom[232][10] = 16'hFFED;
        rom[232][11] = 16'h003E;
        rom[232][12] = 16'hFFD9;
        rom[232][13] = 16'hFFF6;
        rom[232][14] = 16'h0004;
        rom[232][15] = 16'hFFFD;
        rom[232][16] = 16'hFFD7;
        rom[232][17] = 16'hFFCC;
        rom[232][18] = 16'h002A;
        rom[232][19] = 16'hFFDE;
        rom[232][20] = 16'hFFF8;
        rom[232][21] = 16'hFFE8;
        rom[232][22] = 16'h000C;
        rom[232][23] = 16'h0027;
        rom[232][24] = 16'hFFF8;
        rom[232][25] = 16'hFFEA;
        rom[232][26] = 16'h0002;
        rom[232][27] = 16'hFFF5;
        rom[232][28] = 16'h000A;
        rom[232][29] = 16'h000B;
        rom[232][30] = 16'hFFE9;
        rom[232][31] = 16'hFFFC;
        rom[232][32] = 16'h000F;
        rom[232][33] = 16'hFFDC;
        rom[232][34] = 16'hFFFE;
        rom[232][35] = 16'h0006;
        rom[232][36] = 16'hFFDA;
        rom[232][37] = 16'hFFE4;
        rom[232][38] = 16'hFFFA;
        rom[232][39] = 16'hFFEB;
        rom[232][40] = 16'hFFE7;
        rom[232][41] = 16'hFFD2;
        rom[232][42] = 16'hFFEA;
        rom[232][43] = 16'h000C;
        rom[232][44] = 16'hFFC1;
        rom[232][45] = 16'hFFFF;
        rom[232][46] = 16'h0016;
        rom[232][47] = 16'h001F;
        rom[232][48] = 16'hFFD1;
        rom[232][49] = 16'hFFC7;
        rom[232][50] = 16'hFFF1;
        rom[232][51] = 16'hFFEF;
        rom[232][52] = 16'hFFFA;
        rom[232][53] = 16'h0015;
        rom[232][54] = 16'hFFD9;
        rom[232][55] = 16'hFFBF;
        rom[232][56] = 16'h0024;
        rom[232][57] = 16'hFFC4;
        rom[232][58] = 16'hFFEA;
        rom[232][59] = 16'h000D;
        rom[232][60] = 16'h0009;
        rom[232][61] = 16'hFFE5;
        rom[232][62] = 16'h0001;
        rom[232][63] = 16'hFFFF;
        rom[232][64] = 16'h0006;
        rom[232][65] = 16'hFFC3;
        rom[232][66] = 16'hFFE4;
        rom[232][67] = 16'hFFE7;
        rom[232][68] = 16'hFFCB;
        rom[232][69] = 16'hFFF9;
        rom[232][70] = 16'hFFE7;
        rom[232][71] = 16'hFFF4;
        rom[232][72] = 16'h0025;
        rom[232][73] = 16'hFFE7;
        rom[232][74] = 16'h0009;
        rom[232][75] = 16'hFFEA;
        rom[232][76] = 16'h000B;
        rom[232][77] = 16'hFFEA;
        rom[232][78] = 16'h001F;
        rom[232][79] = 16'hFFB9;
        rom[232][80] = 16'h000D;
        rom[232][81] = 16'hFFF8;
        rom[232][82] = 16'hFFF6;
        rom[232][83] = 16'h001E;
        rom[232][84] = 16'hFFEB;
        rom[232][85] = 16'hFFE1;
        rom[232][86] = 16'hFFFF;
        rom[232][87] = 16'h0001;
        rom[232][88] = 16'hFFB7;
        rom[232][89] = 16'hFFEF;
        rom[232][90] = 16'h0000;
        rom[232][91] = 16'h0002;
        rom[232][92] = 16'h0021;
        rom[232][93] = 16'hFFFB;
        rom[232][94] = 16'h001C;
        rom[232][95] = 16'hFFE6;
        rom[232][96] = 16'hFFFB;
        rom[232][97] = 16'h0009;
        rom[232][98] = 16'hFFEC;
        rom[232][99] = 16'h0000;
        rom[232][100] = 16'h0005;
        rom[232][101] = 16'hFFCA;
        rom[232][102] = 16'hFFFC;
        rom[232][103] = 16'h0015;
        rom[232][104] = 16'hFFF4;
        rom[232][105] = 16'hFFEE;
        rom[232][106] = 16'h002A;
        rom[232][107] = 16'h002B;
        rom[232][108] = 16'h000C;
        rom[232][109] = 16'h0020;
        rom[232][110] = 16'h000F;
        rom[232][111] = 16'h0029;
        rom[232][112] = 16'hFFE7;
        rom[232][113] = 16'hFFD1;
        rom[232][114] = 16'h0011;
        rom[232][115] = 16'h0065;
        rom[232][116] = 16'h0017;
        rom[232][117] = 16'hFFD5;
        rom[232][118] = 16'hFFF0;
        rom[232][119] = 16'hFFF5;
        rom[232][120] = 16'h0017;
        rom[232][121] = 16'h0024;
        rom[232][122] = 16'h0017;
        rom[232][123] = 16'h001F;
        rom[232][124] = 16'hFFE1;
        rom[232][125] = 16'hFFE1;
        rom[232][126] = 16'h001D;
        rom[232][127] = 16'h0021;
        rom[233][0] = 16'hFFE2;
        rom[233][1] = 16'hFFEA;
        rom[233][2] = 16'h0003;
        rom[233][3] = 16'hFFF4;
        rom[233][4] = 16'h0017;
        rom[233][5] = 16'h0029;
        rom[233][6] = 16'hFFDC;
        rom[233][7] = 16'h0013;
        rom[233][8] = 16'hFFC4;
        rom[233][9] = 16'hFFFA;
        rom[233][10] = 16'h0003;
        rom[233][11] = 16'hFFCD;
        rom[233][12] = 16'hFFF6;
        rom[233][13] = 16'h0006;
        rom[233][14] = 16'h0004;
        rom[233][15] = 16'hFFEC;
        rom[233][16] = 16'hFFCF;
        rom[233][17] = 16'h000D;
        rom[233][18] = 16'hFFEB;
        rom[233][19] = 16'hFFCF;
        rom[233][20] = 16'hFFCC;
        rom[233][21] = 16'h0000;
        rom[233][22] = 16'hFFD2;
        rom[233][23] = 16'hFFD3;
        rom[233][24] = 16'h000B;
        rom[233][25] = 16'h0008;
        rom[233][26] = 16'hFFD9;
        rom[233][27] = 16'hFFE6;
        rom[233][28] = 16'h002F;
        rom[233][29] = 16'h001F;
        rom[233][30] = 16'hFFE1;
        rom[233][31] = 16'h0001;
        rom[233][32] = 16'hFFAF;
        rom[233][33] = 16'hFFF4;
        rom[233][34] = 16'hFFEE;
        rom[233][35] = 16'h0028;
        rom[233][36] = 16'hFFF6;
        rom[233][37] = 16'hFFE4;
        rom[233][38] = 16'h0001;
        rom[233][39] = 16'hFFDE;
        rom[233][40] = 16'h0027;
        rom[233][41] = 16'hFFEA;
        rom[233][42] = 16'h0003;
        rom[233][43] = 16'h0011;
        rom[233][44] = 16'h0003;
        rom[233][45] = 16'h0024;
        rom[233][46] = 16'h0011;
        rom[233][47] = 16'h001E;
        rom[233][48] = 16'hFFFA;
        rom[233][49] = 16'h0003;
        rom[233][50] = 16'h0000;
        rom[233][51] = 16'h0001;
        rom[233][52] = 16'h0013;
        rom[233][53] = 16'h0016;
        rom[233][54] = 16'hFFEB;
        rom[233][55] = 16'hFFFD;
        rom[233][56] = 16'hFFEF;
        rom[233][57] = 16'hFFE5;
        rom[233][58] = 16'h0013;
        rom[233][59] = 16'hFFEA;
        rom[233][60] = 16'hFFF3;
        rom[233][61] = 16'hFFD0;
        rom[233][62] = 16'hFFFA;
        rom[233][63] = 16'h0003;
        rom[233][64] = 16'hFFE1;
        rom[233][65] = 16'h0002;
        rom[233][66] = 16'h0029;
        rom[233][67] = 16'hFFEF;
        rom[233][68] = 16'h0006;
        rom[233][69] = 16'hFFF9;
        rom[233][70] = 16'hFFEF;
        rom[233][71] = 16'hFFF6;
        rom[233][72] = 16'hFFF0;
        rom[233][73] = 16'h0011;
        rom[233][74] = 16'h0007;
        rom[233][75] = 16'h0019;
        rom[233][76] = 16'h001F;
        rom[233][77] = 16'h0025;
        rom[233][78] = 16'hFFE0;
        rom[233][79] = 16'hFFEE;
        rom[233][80] = 16'hFFFF;
        rom[233][81] = 16'h0000;
        rom[233][82] = 16'h0013;
        rom[233][83] = 16'hFFEA;
        rom[233][84] = 16'hFFE1;
        rom[233][85] = 16'h000A;
        rom[233][86] = 16'hFFF9;
        rom[233][87] = 16'hFFEF;
        rom[233][88] = 16'hFFDB;
        rom[233][89] = 16'hFFFC;
        rom[233][90] = 16'hFFE8;
        rom[233][91] = 16'hFFDC;
        rom[233][92] = 16'hFFE1;
        rom[233][93] = 16'h0016;
        rom[233][94] = 16'h0013;
        rom[233][95] = 16'hFFD2;
        rom[233][96] = 16'hFFEB;
        rom[233][97] = 16'hFFE5;
        rom[233][98] = 16'hFFE0;
        rom[233][99] = 16'hFFFF;
        rom[233][100] = 16'hFFE1;
        rom[233][101] = 16'hFFE7;
        rom[233][102] = 16'h0018;
        rom[233][103] = 16'hFFED;
        rom[233][104] = 16'h0006;
        rom[233][105] = 16'hFFC0;
        rom[233][106] = 16'h0017;
        rom[233][107] = 16'h0011;
        rom[233][108] = 16'hFFEC;
        rom[233][109] = 16'hFFF6;
        rom[233][110] = 16'h0024;
        rom[233][111] = 16'h0011;
        rom[233][112] = 16'hFFFC;
        rom[233][113] = 16'hFFD2;
        rom[233][114] = 16'hFFE0;
        rom[233][115] = 16'hFFD0;
        rom[233][116] = 16'hFFE5;
        rom[233][117] = 16'hFFF6;
        rom[233][118] = 16'h0041;
        rom[233][119] = 16'h0016;
        rom[233][120] = 16'hFFD2;
        rom[233][121] = 16'hFFEF;
        rom[233][122] = 16'hFFF1;
        rom[233][123] = 16'h0014;
        rom[233][124] = 16'hFFF4;
        rom[233][125] = 16'h000D;
        rom[233][126] = 16'hFFF9;
        rom[233][127] = 16'hFFEE;
        rom[234][0] = 16'hFFD6;
        rom[234][1] = 16'h0002;
        rom[234][2] = 16'h0000;
        rom[234][3] = 16'hFFD5;
        rom[234][4] = 16'hFFE6;
        rom[234][5] = 16'hFFE4;
        rom[234][6] = 16'h0035;
        rom[234][7] = 16'h0007;
        rom[234][8] = 16'hFFFB;
        rom[234][9] = 16'hFFF5;
        rom[234][10] = 16'hFFCF;
        rom[234][11] = 16'hFFEF;
        rom[234][12] = 16'hFFF4;
        rom[234][13] = 16'hFFF1;
        rom[234][14] = 16'h0013;
        rom[234][15] = 16'h001D;
        rom[234][16] = 16'hFFF2;
        rom[234][17] = 16'h0007;
        rom[234][18] = 16'hFFFB;
        rom[234][19] = 16'hFFDC;
        rom[234][20] = 16'hFFD9;
        rom[234][21] = 16'h0020;
        rom[234][22] = 16'hFFE0;
        rom[234][23] = 16'hFFD8;
        rom[234][24] = 16'h0006;
        rom[234][25] = 16'h0019;
        rom[234][26] = 16'hFFF9;
        rom[234][27] = 16'hFFF2;
        rom[234][28] = 16'h0008;
        rom[234][29] = 16'h0004;
        rom[234][30] = 16'h0012;
        rom[234][31] = 16'h0022;
        rom[234][32] = 16'hFFE2;
        rom[234][33] = 16'h0008;
        rom[234][34] = 16'h0003;
        rom[234][35] = 16'h0016;
        rom[234][36] = 16'hFFF1;
        rom[234][37] = 16'hFFE1;
        rom[234][38] = 16'hFFD4;
        rom[234][39] = 16'h0029;
        rom[234][40] = 16'h0008;
        rom[234][41] = 16'hFFD1;
        rom[234][42] = 16'hFFFA;
        rom[234][43] = 16'hFFD1;
        rom[234][44] = 16'h001C;
        rom[234][45] = 16'h0027;
        rom[234][46] = 16'hFFF9;
        rom[234][47] = 16'h0008;
        rom[234][48] = 16'hFFF9;
        rom[234][49] = 16'hFFE9;
        rom[234][50] = 16'h0007;
        rom[234][51] = 16'hFFEA;
        rom[234][52] = 16'h001F;
        rom[234][53] = 16'h000A;
        rom[234][54] = 16'h002E;
        rom[234][55] = 16'h0015;
        rom[234][56] = 16'h000E;
        rom[234][57] = 16'hFFF0;
        rom[234][58] = 16'h000C;
        rom[234][59] = 16'hFFB2;
        rom[234][60] = 16'h0003;
        rom[234][61] = 16'hFFF5;
        rom[234][62] = 16'h0029;
        rom[234][63] = 16'hFFF6;
        rom[234][64] = 16'hFFA0;
        rom[234][65] = 16'h0011;
        rom[234][66] = 16'h000F;
        rom[234][67] = 16'hFFD7;
        rom[234][68] = 16'h0017;
        rom[234][69] = 16'hFFEF;
        rom[234][70] = 16'h002E;
        rom[234][71] = 16'hFFF4;
        rom[234][72] = 16'hFFFB;
        rom[234][73] = 16'h0001;
        rom[234][74] = 16'h000C;
        rom[234][75] = 16'h000F;
        rom[234][76] = 16'hFFF9;
        rom[234][77] = 16'hFFF4;
        rom[234][78] = 16'h000C;
        rom[234][79] = 16'h0016;
        rom[234][80] = 16'h0001;
        rom[234][81] = 16'h001F;
        rom[234][82] = 16'hFFCA;
        rom[234][83] = 16'h0007;
        rom[234][84] = 16'h0007;
        rom[234][85] = 16'h000F;
        rom[234][86] = 16'hFFDE;
        rom[234][87] = 16'h000C;
        rom[234][88] = 16'h000C;
        rom[234][89] = 16'h001F;
        rom[234][90] = 16'hFFBE;
        rom[234][91] = 16'hFFFB;
        rom[234][92] = 16'h001C;
        rom[234][93] = 16'hFFDE;
        rom[234][94] = 16'hFFF5;
        rom[234][95] = 16'hFFBF;
        rom[234][96] = 16'hFFFC;
        rom[234][97] = 16'hFFF7;
        rom[234][98] = 16'hFFF9;
        rom[234][99] = 16'h0002;
        rom[234][100] = 16'h0005;
        rom[234][101] = 16'hFFB0;
        rom[234][102] = 16'hFFF7;
        rom[234][103] = 16'h0066;
        rom[234][104] = 16'hFFD4;
        rom[234][105] = 16'h0015;
        rom[234][106] = 16'hFFE0;
        rom[234][107] = 16'h000C;
        rom[234][108] = 16'h0002;
        rom[234][109] = 16'hFFCD;
        rom[234][110] = 16'hFFEF;
        rom[234][111] = 16'hFFEC;
        rom[234][112] = 16'hFFE1;
        rom[234][113] = 16'h0007;
        rom[234][114] = 16'h0003;
        rom[234][115] = 16'h0045;
        rom[234][116] = 16'h0016;
        rom[234][117] = 16'hFFD3;
        rom[234][118] = 16'hFFDB;
        rom[234][119] = 16'h001E;
        rom[234][120] = 16'h000D;
        rom[234][121] = 16'hFFCF;
        rom[234][122] = 16'h0015;
        rom[234][123] = 16'hFFFE;
        rom[234][124] = 16'h002C;
        rom[234][125] = 16'h0015;
        rom[234][126] = 16'h000C;
        rom[234][127] = 16'hFFF1;
        rom[235][0] = 16'hFFF9;
        rom[235][1] = 16'hFFF4;
        rom[235][2] = 16'h0039;
        rom[235][3] = 16'h0011;
        rom[235][4] = 16'h000C;
        rom[235][5] = 16'h0003;
        rom[235][6] = 16'hFFF3;
        rom[235][7] = 16'h001B;
        rom[235][8] = 16'h0043;
        rom[235][9] = 16'h0019;
        rom[235][10] = 16'h0007;
        rom[235][11] = 16'h0002;
        rom[235][12] = 16'hFFEA;
        rom[235][13] = 16'hFFE7;
        rom[235][14] = 16'h0020;
        rom[235][15] = 16'hFFFD;
        rom[235][16] = 16'hFFCA;
        rom[235][17] = 16'hFFDB;
        rom[235][18] = 16'h0016;
        rom[235][19] = 16'h000C;
        rom[235][20] = 16'h0029;
        rom[235][21] = 16'h0025;
        rom[235][22] = 16'hFFE5;
        rom[235][23] = 16'h0007;
        rom[235][24] = 16'hFFEF;
        rom[235][25] = 16'h004E;
        rom[235][26] = 16'h002E;
        rom[235][27] = 16'hFFDA;
        rom[235][28] = 16'hFFEE;
        rom[235][29] = 16'h001B;
        rom[235][30] = 16'h0024;
        rom[235][31] = 16'h0037;
        rom[235][32] = 16'h003F;
        rom[235][33] = 16'hFFD0;
        rom[235][34] = 16'h0002;
        rom[235][35] = 16'hFFD2;
        rom[235][36] = 16'h0036;
        rom[235][37] = 16'h0007;
        rom[235][38] = 16'h0004;
        rom[235][39] = 16'hFFB5;
        rom[235][40] = 16'h0000;
        rom[235][41] = 16'h0015;
        rom[235][42] = 16'h0014;
        rom[235][43] = 16'hFFEC;
        rom[235][44] = 16'hFFFB;
        rom[235][45] = 16'hFFE9;
        rom[235][46] = 16'hFFE5;
        rom[235][47] = 16'h000A;
        rom[235][48] = 16'h0012;
        rom[235][49] = 16'h000C;
        rom[235][50] = 16'hFFD1;
        rom[235][51] = 16'hFFFE;
        rom[235][52] = 16'hFFC5;
        rom[235][53] = 16'h0011;
        rom[235][54] = 16'hFFEB;
        rom[235][55] = 16'h0055;
        rom[235][56] = 16'h0028;
        rom[235][57] = 16'hFFB3;
        rom[235][58] = 16'hFFE3;
        rom[235][59] = 16'h001A;
        rom[235][60] = 16'hFFF7;
        rom[235][61] = 16'h0005;
        rom[235][62] = 16'hFFDA;
        rom[235][63] = 16'hFFFE;
        rom[235][64] = 16'h000E;
        rom[235][65] = 16'h0013;
        rom[235][66] = 16'h0000;
        rom[235][67] = 16'hFFFE;
        rom[235][68] = 16'h001D;
        rom[235][69] = 16'h0001;
        rom[235][70] = 16'h001B;
        rom[235][71] = 16'h0028;
        rom[235][72] = 16'h001C;
        rom[235][73] = 16'hFFF1;
        rom[235][74] = 16'h0034;
        rom[235][75] = 16'hFFD5;
        rom[235][76] = 16'hFFFE;
        rom[235][77] = 16'hFFCA;
        rom[235][78] = 16'h0007;
        rom[235][79] = 16'h0004;
        rom[235][80] = 16'h0003;
        rom[235][81] = 16'hFFCF;
        rom[235][82] = 16'h0015;
        rom[235][83] = 16'h003E;
        rom[235][84] = 16'h0033;
        rom[235][85] = 16'hFFDB;
        rom[235][86] = 16'hFFF3;
        rom[235][87] = 16'hFFC7;
        rom[235][88] = 16'hFFFD;
        rom[235][89] = 16'hFFC3;
        rom[235][90] = 16'h002F;
        rom[235][91] = 16'hFFDB;
        rom[235][92] = 16'hFFDD;
        rom[235][93] = 16'hFFB0;
        rom[235][94] = 16'h0004;
        rom[235][95] = 16'hFFEB;
        rom[235][96] = 16'hFFC1;
        rom[235][97] = 16'h0004;
        rom[235][98] = 16'hFFCF;
        rom[235][99] = 16'hFFF0;
        rom[235][100] = 16'hFFDA;
        rom[235][101] = 16'h0044;
        rom[235][102] = 16'hFFE2;
        rom[235][103] = 16'hFFDA;
        rom[235][104] = 16'h002E;
        rom[235][105] = 16'h0044;
        rom[235][106] = 16'h000E;
        rom[235][107] = 16'hFFF1;
        rom[235][108] = 16'h002D;
        rom[235][109] = 16'hFFEC;
        rom[235][110] = 16'h002F;
        rom[235][111] = 16'hFFFB;
        rom[235][112] = 16'h0011;
        rom[235][113] = 16'h001B;
        rom[235][114] = 16'hFFEA;
        rom[235][115] = 16'h0016;
        rom[235][116] = 16'hFFB0;
        rom[235][117] = 16'hFFF6;
        rom[235][118] = 16'hFFF0;
        rom[235][119] = 16'hFFEF;
        rom[235][120] = 16'h000D;
        rom[235][121] = 16'hFFD4;
        rom[235][122] = 16'hFFF2;
        rom[235][123] = 16'hFFB3;
        rom[235][124] = 16'hFFBE;
        rom[235][125] = 16'h0002;
        rom[235][126] = 16'hFFDE;
        rom[235][127] = 16'hFFF2;
        rom[236][0] = 16'hFFC3;
        rom[236][1] = 16'h0015;
        rom[236][2] = 16'h0011;
        rom[236][3] = 16'hFFCD;
        rom[236][4] = 16'hFFD7;
        rom[236][5] = 16'h0006;
        rom[236][6] = 16'h0014;
        rom[236][7] = 16'hFFEE;
        rom[236][8] = 16'h001D;
        rom[236][9] = 16'hFFEA;
        rom[236][10] = 16'h0012;
        rom[236][11] = 16'hFFD7;
        rom[236][12] = 16'h0005;
        rom[236][13] = 16'h0012;
        rom[236][14] = 16'h0002;
        rom[236][15] = 16'h0001;
        rom[236][16] = 16'h0008;
        rom[236][17] = 16'hFFDC;
        rom[236][18] = 16'hFFD0;
        rom[236][19] = 16'h0020;
        rom[236][20] = 16'h000D;
        rom[236][21] = 16'h0017;
        rom[236][22] = 16'hFFFC;
        rom[236][23] = 16'hFFDF;
        rom[236][24] = 16'hFFFB;
        rom[236][25] = 16'h0036;
        rom[236][26] = 16'hFFC2;
        rom[236][27] = 16'h0036;
        rom[236][28] = 16'h0005;
        rom[236][29] = 16'h0010;
        rom[236][30] = 16'h0008;
        rom[236][31] = 16'h001B;
        rom[236][32] = 16'hFFD4;
        rom[236][33] = 16'hFFEE;
        rom[236][34] = 16'h001A;
        rom[236][35] = 16'h001B;
        rom[236][36] = 16'h0006;
        rom[236][37] = 16'hFFAC;
        rom[236][38] = 16'hFFD1;
        rom[236][39] = 16'hFFF8;
        rom[236][40] = 16'h0022;
        rom[236][41] = 16'hFFF4;
        rom[236][42] = 16'h003B;
        rom[236][43] = 16'hFFE0;
        rom[236][44] = 16'h0006;
        rom[236][45] = 16'h0027;
        rom[236][46] = 16'h0012;
        rom[236][47] = 16'h0029;
        rom[236][48] = 16'hFFF9;
        rom[236][49] = 16'h0029;
        rom[236][50] = 16'h0004;
        rom[236][51] = 16'hFFBA;
        rom[236][52] = 16'hFFDD;
        rom[236][53] = 16'h0011;
        rom[236][54] = 16'hFFFE;
        rom[236][55] = 16'h001B;
        rom[236][56] = 16'h000E;
        rom[236][57] = 16'hFFDC;
        rom[236][58] = 16'hFFFF;
        rom[236][59] = 16'hFFDC;
        rom[236][60] = 16'h001F;
        rom[236][61] = 16'h0007;
        rom[236][62] = 16'h002C;
        rom[236][63] = 16'h0001;
        rom[236][64] = 16'hFFC3;
        rom[236][65] = 16'h000F;
        rom[236][66] = 16'hFFF1;
        rom[236][67] = 16'h0009;
        rom[236][68] = 16'hFFD2;
        rom[236][69] = 16'hFFFF;
        rom[236][70] = 16'h0020;
        rom[236][71] = 16'hFFCC;
        rom[236][72] = 16'h0002;
        rom[236][73] = 16'hFFFE;
        rom[236][74] = 16'hFFE6;
        rom[236][75] = 16'hFFE3;
        rom[236][76] = 16'h0016;
        rom[236][77] = 16'hFFD7;
        rom[236][78] = 16'hFFFB;
        rom[236][79] = 16'h0007;
        rom[236][80] = 16'h0009;
        rom[236][81] = 16'h0011;
        rom[236][82] = 16'hFFF4;
        rom[236][83] = 16'h0011;
        rom[236][84] = 16'h0005;
        rom[236][85] = 16'hFFDF;
        rom[236][86] = 16'hFFE9;
        rom[236][87] = 16'hFFDA;
        rom[236][88] = 16'h0013;
        rom[236][89] = 16'h0013;
        rom[236][90] = 16'h0001;
        rom[236][91] = 16'hFFEF;
        rom[236][92] = 16'hFFFE;
        rom[236][93] = 16'hFFF0;
        rom[236][94] = 16'hFF9F;
        rom[236][95] = 16'hFFBA;
        rom[236][96] = 16'h0016;
        rom[236][97] = 16'hFFF4;
        rom[236][98] = 16'h0014;
        rom[236][99] = 16'h0024;
        rom[236][100] = 16'h001B;
        rom[236][101] = 16'hFFE3;
        rom[236][102] = 16'hFFF9;
        rom[236][103] = 16'hFFD5;
        rom[236][104] = 16'hFFD6;
        rom[236][105] = 16'hFFB9;
        rom[236][106] = 16'h0005;
        rom[236][107] = 16'h000E;
        rom[236][108] = 16'h0001;
        rom[236][109] = 16'hFFE5;
        rom[236][110] = 16'h0000;
        rom[236][111] = 16'h0000;
        rom[236][112] = 16'hFFD9;
        rom[236][113] = 16'h0011;
        rom[236][114] = 16'h0019;
        rom[236][115] = 16'h0034;
        rom[236][116] = 16'hFFC8;
        rom[236][117] = 16'hFFD2;
        rom[236][118] = 16'hFFFB;
        rom[236][119] = 16'h0039;
        rom[236][120] = 16'hFFF2;
        rom[236][121] = 16'hFFF3;
        rom[236][122] = 16'hFFFF;
        rom[236][123] = 16'hFFE5;
        rom[236][124] = 16'hFFEF;
        rom[236][125] = 16'hFFBC;
        rom[236][126] = 16'h0011;
        rom[236][127] = 16'hFFD8;
        rom[237][0] = 16'h0009;
        rom[237][1] = 16'h0021;
        rom[237][2] = 16'hFFDD;
        rom[237][3] = 16'hFFE9;
        rom[237][4] = 16'hFFFD;
        rom[237][5] = 16'hFFEB;
        rom[237][6] = 16'hFFFA;
        rom[237][7] = 16'hFFCA;
        rom[237][8] = 16'h0010;
        rom[237][9] = 16'hFFE1;
        rom[237][10] = 16'hFFF0;
        rom[237][11] = 16'h0020;
        rom[237][12] = 16'hFFF7;
        rom[237][13] = 16'hFFE6;
        rom[237][14] = 16'h000C;
        rom[237][15] = 16'h0008;
        rom[237][16] = 16'h0003;
        rom[237][17] = 16'hFFB6;
        rom[237][18] = 16'hFFCB;
        rom[237][19] = 16'h0011;
        rom[237][20] = 16'h001E;
        rom[237][21] = 16'hFFD3;
        rom[237][22] = 16'hFFD0;
        rom[237][23] = 16'h0012;
        rom[237][24] = 16'h0018;
        rom[237][25] = 16'h000E;
        rom[237][26] = 16'h000B;
        rom[237][27] = 16'h0020;
        rom[237][28] = 16'h0016;
        rom[237][29] = 16'h001B;
        rom[237][30] = 16'hFFD6;
        rom[237][31] = 16'h0016;
        rom[237][32] = 16'hFFF3;
        rom[237][33] = 16'hFFAB;
        rom[237][34] = 16'hFFF7;
        rom[237][35] = 16'h002C;
        rom[237][36] = 16'hFFF4;
        rom[237][37] = 16'hFFF4;
        rom[237][38] = 16'hFF9B;
        rom[237][39] = 16'h0031;
        rom[237][40] = 16'hFF9F;
        rom[237][41] = 16'h000F;
        rom[237][42] = 16'hFFF1;
        rom[237][43] = 16'hFFD3;
        rom[237][44] = 16'h0010;
        rom[237][45] = 16'hFFFC;
        rom[237][46] = 16'h000F;
        rom[237][47] = 16'h0007;
        rom[237][48] = 16'hFFDE;
        rom[237][49] = 16'hFFE5;
        rom[237][50] = 16'hFFBB;
        rom[237][51] = 16'hFFDA;
        rom[237][52] = 16'h0003;
        rom[237][53] = 16'hFFEF;
        rom[237][54] = 16'h0001;
        rom[237][55] = 16'h0028;
        rom[237][56] = 16'hFFC0;
        rom[237][57] = 16'hFFFD;
        rom[237][58] = 16'h0016;
        rom[237][59] = 16'h0017;
        rom[237][60] = 16'hFFF4;
        rom[237][61] = 16'h001F;
        rom[237][62] = 16'h0007;
        rom[237][63] = 16'hFFE7;
        rom[237][64] = 16'h0000;
        rom[237][65] = 16'hFFC3;
        rom[237][66] = 16'h0012;
        rom[237][67] = 16'hFFE3;
        rom[237][68] = 16'hFFD0;
        rom[237][69] = 16'h0022;
        rom[237][70] = 16'hFFC3;
        rom[237][71] = 16'hFFF1;
        rom[237][72] = 16'hFFEF;
        rom[237][73] = 16'hFFE7;
        rom[237][74] = 16'hFFC6;
        rom[237][75] = 16'hFFB9;
        rom[237][76] = 16'hFFFB;
        rom[237][77] = 16'hFFF1;
        rom[237][78] = 16'h0007;
        rom[237][79] = 16'h0018;
        rom[237][80] = 16'h0012;
        rom[237][81] = 16'hFFF4;
        rom[237][82] = 16'h0003;
        rom[237][83] = 16'h0018;
        rom[237][84] = 16'h0016;
        rom[237][85] = 16'hFFDF;
        rom[237][86] = 16'hFFFF;
        rom[237][87] = 16'hFFF5;
        rom[237][88] = 16'hFFDA;
        rom[237][89] = 16'hFFF5;
        rom[237][90] = 16'h000C;
        rom[237][91] = 16'hFFEA;
        rom[237][92] = 16'hFFD9;
        rom[237][93] = 16'h0006;
        rom[237][94] = 16'hFFA2;
        rom[237][95] = 16'h000A;
        rom[237][96] = 16'hFFEB;
        rom[237][97] = 16'h000D;
        rom[237][98] = 16'h0004;
        rom[237][99] = 16'h001B;
        rom[237][100] = 16'h0006;
        rom[237][101] = 16'h000C;
        rom[237][102] = 16'hFFE2;
        rom[237][103] = 16'hFFFA;
        rom[237][104] = 16'hFFD7;
        rom[237][105] = 16'h0030;
        rom[237][106] = 16'hFFD9;
        rom[237][107] = 16'h0016;
        rom[237][108] = 16'h0008;
        rom[237][109] = 16'hFFEA;
        rom[237][110] = 16'h0017;
        rom[237][111] = 16'h000C;
        rom[237][112] = 16'h0012;
        rom[237][113] = 16'h0013;
        rom[237][114] = 16'hFFF1;
        rom[237][115] = 16'hFFE8;
        rom[237][116] = 16'h000F;
        rom[237][117] = 16'h000B;
        rom[237][118] = 16'h0014;
        rom[237][119] = 16'hFFE4;
        rom[237][120] = 16'hFFCD;
        rom[237][121] = 16'h000C;
        rom[237][122] = 16'hFFE7;
        rom[237][123] = 16'hFFC5;
        rom[237][124] = 16'hFFFE;
        rom[237][125] = 16'hFFE4;
        rom[237][126] = 16'hFFEB;
        rom[237][127] = 16'hFFFE;
        rom[238][0] = 16'h0016;
        rom[238][1] = 16'hFFB0;
        rom[238][2] = 16'hFFEF;
        rom[238][3] = 16'h0015;
        rom[238][4] = 16'hFFC3;
        rom[238][5] = 16'hFFDC;
        rom[238][6] = 16'h0006;
        rom[238][7] = 16'hFFFF;
        rom[238][8] = 16'hFFFA;
        rom[238][9] = 16'h001F;
        rom[238][10] = 16'h0025;
        rom[238][11] = 16'h0017;
        rom[238][12] = 16'hFFF1;
        rom[238][13] = 16'h0016;
        rom[238][14] = 16'h0007;
        rom[238][15] = 16'h0001;
        rom[238][16] = 16'h000F;
        rom[238][17] = 16'h0022;
        rom[238][18] = 16'hFFF3;
        rom[238][19] = 16'h0003;
        rom[238][20] = 16'hFFF4;
        rom[238][21] = 16'hFFC1;
        rom[238][22] = 16'h0016;
        rom[238][23] = 16'h0014;
        rom[238][24] = 16'h001B;
        rom[238][25] = 16'hFFDF;
        rom[238][26] = 16'h0006;
        rom[238][27] = 16'hFFD9;
        rom[238][28] = 16'hFFB7;
        rom[238][29] = 16'h000F;
        rom[238][30] = 16'hFFEA;
        rom[238][31] = 16'hFFFC;
        rom[238][32] = 16'hFFFA;
        rom[238][33] = 16'h0020;
        rom[238][34] = 16'h000A;
        rom[238][35] = 16'h0003;
        rom[238][36] = 16'hFFEE;
        rom[238][37] = 16'hFFB8;
        rom[238][38] = 16'h0000;
        rom[238][39] = 16'h001A;
        rom[238][40] = 16'h0015;
        rom[238][41] = 16'h000C;
        rom[238][42] = 16'hFFD6;
        rom[238][43] = 16'h0003;
        rom[238][44] = 16'h0029;
        rom[238][45] = 16'hFFF7;
        rom[238][46] = 16'hFFD8;
        rom[238][47] = 16'hFFFF;
        rom[238][48] = 16'h0022;
        rom[238][49] = 16'hFFFB;
        rom[238][50] = 16'h000A;
        rom[238][51] = 16'hFFFE;
        rom[238][52] = 16'hFFDF;
        rom[238][53] = 16'h003A;
        rom[238][54] = 16'hFFC2;
        rom[238][55] = 16'hFFFD;
        rom[238][56] = 16'h0000;
        rom[238][57] = 16'h001D;
        rom[238][58] = 16'hFFDE;
        rom[238][59] = 16'hFFFD;
        rom[238][60] = 16'hFFE1;
        rom[238][61] = 16'hFFD3;
        rom[238][62] = 16'hFFE3;
        rom[238][63] = 16'hFFED;
        rom[238][64] = 16'hFFD4;
        rom[238][65] = 16'hFFDA;
        rom[238][66] = 16'hFFEB;
        rom[238][67] = 16'hFFED;
        rom[238][68] = 16'h001E;
        rom[238][69] = 16'hFFDA;
        rom[238][70] = 16'hFFDF;
        rom[238][71] = 16'hFFAC;
        rom[238][72] = 16'hFFE5;
        rom[238][73] = 16'h001F;
        rom[238][74] = 16'h000F;
        rom[238][75] = 16'hFFF9;
        rom[238][76] = 16'hFFF8;
        rom[238][77] = 16'h0017;
        rom[238][78] = 16'h0008;
        rom[238][79] = 16'hFFD5;
        rom[238][80] = 16'hFFEE;
        rom[238][81] = 16'hFFF4;
        rom[238][82] = 16'hFFAB;
        rom[238][83] = 16'h0006;
        rom[238][84] = 16'hFFFF;
        rom[238][85] = 16'hFFD5;
        rom[238][86] = 16'hFFF4;
        rom[238][87] = 16'h0014;
        rom[238][88] = 16'h0008;
        rom[238][89] = 16'hFFF4;
        rom[238][90] = 16'hFFD9;
        rom[238][91] = 16'h000D;
        rom[238][92] = 16'hFFF2;
        rom[238][93] = 16'h0025;
        rom[238][94] = 16'h002D;
        rom[238][95] = 16'hFFEC;
        rom[238][96] = 16'h0005;
        rom[238][97] = 16'h0031;
        rom[238][98] = 16'hFFF6;
        rom[238][99] = 16'hFFF3;
        rom[238][100] = 16'hFFFF;
        rom[238][101] = 16'h0010;
        rom[238][102] = 16'h0006;
        rom[238][103] = 16'h001E;
        rom[238][104] = 16'hFFFC;
        rom[238][105] = 16'hFFF4;
        rom[238][106] = 16'h0000;
        rom[238][107] = 16'h0002;
        rom[238][108] = 16'hFFE0;
        rom[238][109] = 16'hFFDA;
        rom[238][110] = 16'hFFD2;
        rom[238][111] = 16'h0001;
        rom[238][112] = 16'hFFCF;
        rom[238][113] = 16'hFFEA;
        rom[238][114] = 16'h0002;
        rom[238][115] = 16'h0017;
        rom[238][116] = 16'hFFCD;
        rom[238][117] = 16'hFFF5;
        rom[238][118] = 16'hFFD2;
        rom[238][119] = 16'hFFFD;
        rom[238][120] = 16'h0006;
        rom[238][121] = 16'h0002;
        rom[238][122] = 16'hFFFF;
        rom[238][123] = 16'hFFE3;
        rom[238][124] = 16'hFFF1;
        rom[238][125] = 16'hFFFB;
        rom[238][126] = 16'hFFE0;
        rom[238][127] = 16'h002D;
        rom[239][0] = 16'hFFF1;
        rom[239][1] = 16'h0007;
        rom[239][2] = 16'h0011;
        rom[239][3] = 16'h0005;
        rom[239][4] = 16'hFFFC;
        rom[239][5] = 16'hFFD6;
        rom[239][6] = 16'h002B;
        rom[239][7] = 16'h0007;
        rom[239][8] = 16'hFFE8;
        rom[239][9] = 16'h0016;
        rom[239][10] = 16'hFFD9;
        rom[239][11] = 16'h0023;
        rom[239][12] = 16'hFFE2;
        rom[239][13] = 16'h0021;
        rom[239][14] = 16'h0016;
        rom[239][15] = 16'hFFF2;
        rom[239][16] = 16'h0021;
        rom[239][17] = 16'h0001;
        rom[239][18] = 16'h0037;
        rom[239][19] = 16'h001C;
        rom[239][20] = 16'h002D;
        rom[239][21] = 16'hFFB8;
        rom[239][22] = 16'hFFF7;
        rom[239][23] = 16'hFFE1;
        rom[239][24] = 16'h000E;
        rom[239][25] = 16'h0007;
        rom[239][26] = 16'hFFE9;
        rom[239][27] = 16'hFFE2;
        rom[239][28] = 16'hFFE2;
        rom[239][29] = 16'h0019;
        rom[239][30] = 16'h0000;
        rom[239][31] = 16'hFFFC;
        rom[239][32] = 16'h0011;
        rom[239][33] = 16'h001A;
        rom[239][34] = 16'h0002;
        rom[239][35] = 16'hFFE4;
        rom[239][36] = 16'h0038;
        rom[239][37] = 16'hFFDE;
        rom[239][38] = 16'hFFF1;
        rom[239][39] = 16'hFFF1;
        rom[239][40] = 16'h0021;
        rom[239][41] = 16'hFFD2;
        rom[239][42] = 16'h0028;
        rom[239][43] = 16'h0002;
        rom[239][44] = 16'h0007;
        rom[239][45] = 16'hFFF2;
        rom[239][46] = 16'h0030;
        rom[239][47] = 16'hFFF5;
        rom[239][48] = 16'h000B;
        rom[239][49] = 16'h0037;
        rom[239][50] = 16'hFFEF;
        rom[239][51] = 16'h001B;
        rom[239][52] = 16'hFFD7;
        rom[239][53] = 16'h0028;
        rom[239][54] = 16'hFFFE;
        rom[239][55] = 16'h0068;
        rom[239][56] = 16'h0014;
        rom[239][57] = 16'h0030;
        rom[239][58] = 16'h0026;
        rom[239][59] = 16'hFFD0;
        rom[239][60] = 16'hFFD1;
        rom[239][61] = 16'h001A;
        rom[239][62] = 16'h0022;
        rom[239][63] = 16'hFFF9;
        rom[239][64] = 16'h0033;
        rom[239][65] = 16'h002A;
        rom[239][66] = 16'hFFC2;
        rom[239][67] = 16'hFFD1;
        rom[239][68] = 16'h0039;
        rom[239][69] = 16'hFFD2;
        rom[239][70] = 16'hFFE1;
        rom[239][71] = 16'h0006;
        rom[239][72] = 16'h0015;
        rom[239][73] = 16'hFFF1;
        rom[239][74] = 16'hFFF7;
        rom[239][75] = 16'hFFFF;
        rom[239][76] = 16'h0004;
        rom[239][77] = 16'h0007;
        rom[239][78] = 16'hFFFE;
        rom[239][79] = 16'h0009;
        rom[239][80] = 16'h000A;
        rom[239][81] = 16'h000B;
        rom[239][82] = 16'hFFF9;
        rom[239][83] = 16'hFFAE;
        rom[239][84] = 16'h0023;
        rom[239][85] = 16'h001A;
        rom[239][86] = 16'h002D;
        rom[239][87] = 16'hFFE7;
        rom[239][88] = 16'hFFE3;
        rom[239][89] = 16'hFFE5;
        rom[239][90] = 16'h0003;
        rom[239][91] = 16'hFFF9;
        rom[239][92] = 16'hFFDF;
        rom[239][93] = 16'hFFED;
        rom[239][94] = 16'h0037;
        rom[239][95] = 16'hFFBF;
        rom[239][96] = 16'h0009;
        rom[239][97] = 16'hFFFA;
        rom[239][98] = 16'hFFEF;
        rom[239][99] = 16'hFFF4;
        rom[239][100] = 16'hFFEF;
        rom[239][101] = 16'hFFCD;
        rom[239][102] = 16'h0014;
        rom[239][103] = 16'hFFF7;
        rom[239][104] = 16'h000C;
        rom[239][105] = 16'hFFD2;
        rom[239][106] = 16'h0006;
        rom[239][107] = 16'hFFE0;
        rom[239][108] = 16'h000C;
        rom[239][109] = 16'hFFCC;
        rom[239][110] = 16'h0001;
        rom[239][111] = 16'hFFBA;
        rom[239][112] = 16'hFFF8;
        rom[239][113] = 16'h0015;
        rom[239][114] = 16'hFFF7;
        rom[239][115] = 16'h0012;
        rom[239][116] = 16'h0025;
        rom[239][117] = 16'hFFF0;
        rom[239][118] = 16'hFFEA;
        rom[239][119] = 16'h001C;
        rom[239][120] = 16'h0024;
        rom[239][121] = 16'h000A;
        rom[239][122] = 16'hFFF7;
        rom[239][123] = 16'hFFF6;
        rom[239][124] = 16'h001C;
        rom[239][125] = 16'hFFF7;
        rom[239][126] = 16'hFFDD;
        rom[239][127] = 16'hFFD1;
        rom[240][0] = 16'hFFD4;
        rom[240][1] = 16'h0019;
        rom[240][2] = 16'hFFD2;
        rom[240][3] = 16'hFFC0;
        rom[240][4] = 16'hFFEF;
        rom[240][5] = 16'hFFDB;
        rom[240][6] = 16'h000C;
        rom[240][7] = 16'hFFEF;
        rom[240][8] = 16'h001F;
        rom[240][9] = 16'hFFD9;
        rom[240][10] = 16'hFFD7;
        rom[240][11] = 16'h0005;
        rom[240][12] = 16'h0021;
        rom[240][13] = 16'h0011;
        rom[240][14] = 16'h0011;
        rom[240][15] = 16'h001C;
        rom[240][16] = 16'hFFFE;
        rom[240][17] = 16'h0007;
        rom[240][18] = 16'hFFAC;
        rom[240][19] = 16'h0007;
        rom[240][20] = 16'hFFDA;
        rom[240][21] = 16'hFFC5;
        rom[240][22] = 16'hFFE7;
        rom[240][23] = 16'hFFB7;
        rom[240][24] = 16'h001B;
        rom[240][25] = 16'h0000;
        rom[240][26] = 16'hFFEF;
        rom[240][27] = 16'hFFFE;
        rom[240][28] = 16'h0011;
        rom[240][29] = 16'h0017;
        rom[240][30] = 16'hFFFE;
        rom[240][31] = 16'h000A;
        rom[240][32] = 16'h0018;
        rom[240][33] = 16'h0008;
        rom[240][34] = 16'hFFE1;
        rom[240][35] = 16'hFFF9;
        rom[240][36] = 16'hFFF7;
        rom[240][37] = 16'h0016;
        rom[240][38] = 16'hFFFE;
        rom[240][39] = 16'h000D;
        rom[240][40] = 16'hFFF8;
        rom[240][41] = 16'h001B;
        rom[240][42] = 16'hFFFB;
        rom[240][43] = 16'hFFE4;
        rom[240][44] = 16'hFFF3;
        rom[240][45] = 16'h000D;
        rom[240][46] = 16'hFFD5;
        rom[240][47] = 16'hFFEA;
        rom[240][48] = 16'h0011;
        rom[240][49] = 16'h0008;
        rom[240][50] = 16'hFFF6;
        rom[240][51] = 16'h0011;
        rom[240][52] = 16'hFFEB;
        rom[240][53] = 16'hFFFD;
        rom[240][54] = 16'h0000;
        rom[240][55] = 16'hFFED;
        rom[240][56] = 16'h000F;
        rom[240][57] = 16'hFFFE;
        rom[240][58] = 16'h0014;
        rom[240][59] = 16'hFFF4;
        rom[240][60] = 16'hFFDD;
        rom[240][61] = 16'h0007;
        rom[240][62] = 16'h003A;
        rom[240][63] = 16'h000E;
        rom[240][64] = 16'h0036;
        rom[240][65] = 16'h0013;
        rom[240][66] = 16'hFFF6;
        rom[240][67] = 16'h0006;
        rom[240][68] = 16'h0009;
        rom[240][69] = 16'h0005;
        rom[240][70] = 16'h0006;
        rom[240][71] = 16'hFFCC;
        rom[240][72] = 16'hFFF4;
        rom[240][73] = 16'h0031;
        rom[240][74] = 16'h0001;
        rom[240][75] = 16'h0004;
        rom[240][76] = 16'hFFEE;
        rom[240][77] = 16'hFFF7;
        rom[240][78] = 16'h002C;
        rom[240][79] = 16'h0045;
        rom[240][80] = 16'hFFE8;
        rom[240][81] = 16'h0009;
        rom[240][82] = 16'h000F;
        rom[240][83] = 16'h0000;
        rom[240][84] = 16'h002B;
        rom[240][85] = 16'h0002;
        rom[240][86] = 16'hFFBF;
        rom[240][87] = 16'h0021;
        rom[240][88] = 16'h0009;
        rom[240][89] = 16'h0015;
        rom[240][90] = 16'hFFF0;
        rom[240][91] = 16'hFFE4;
        rom[240][92] = 16'h000D;
        rom[240][93] = 16'hFFED;
        rom[240][94] = 16'h0005;
        rom[240][95] = 16'h003C;
        rom[240][96] = 16'h0015;
        rom[240][97] = 16'h0021;
        rom[240][98] = 16'hFFBA;
        rom[240][99] = 16'h0003;
        rom[240][100] = 16'hFFEA;
        rom[240][101] = 16'hFFC1;
        rom[240][102] = 16'hFFEA;
        rom[240][103] = 16'hFFD0;
        rom[240][104] = 16'h0002;
        rom[240][105] = 16'hFFF9;
        rom[240][106] = 16'hFFFF;
        rom[240][107] = 16'hFFE5;
        rom[240][108] = 16'hFFEC;
        rom[240][109] = 16'h0033;
        rom[240][110] = 16'h0017;
        rom[240][111] = 16'hFFCF;
        rom[240][112] = 16'h0001;
        rom[240][113] = 16'h001C;
        rom[240][114] = 16'hFFCC;
        rom[240][115] = 16'h0007;
        rom[240][116] = 16'h000C;
        rom[240][117] = 16'hFFF9;
        rom[240][118] = 16'hFFD5;
        rom[240][119] = 16'h0026;
        rom[240][120] = 16'h0002;
        rom[240][121] = 16'hFFB8;
        rom[240][122] = 16'h0011;
        rom[240][123] = 16'hFFED;
        rom[240][124] = 16'h0029;
        rom[240][125] = 16'h0013;
        rom[240][126] = 16'hFFF0;
        rom[240][127] = 16'hFFBF;
        rom[241][0] = 16'hFFD3;
        rom[241][1] = 16'h0029;
        rom[241][2] = 16'h0002;
        rom[241][3] = 16'h002E;
        rom[241][4] = 16'hFFF4;
        rom[241][5] = 16'h0018;
        rom[241][6] = 16'hFFE0;
        rom[241][7] = 16'hFFFC;
        rom[241][8] = 16'hFFFE;
        rom[241][9] = 16'h0008;
        rom[241][10] = 16'h000B;
        rom[241][11] = 16'hFFED;
        rom[241][12] = 16'hFFC7;
        rom[241][13] = 16'h0007;
        rom[241][14] = 16'hFFD8;
        rom[241][15] = 16'h0014;
        rom[241][16] = 16'h0009;
        rom[241][17] = 16'h0016;
        rom[241][18] = 16'hFFE5;
        rom[241][19] = 16'hFFFD;
        rom[241][20] = 16'hFFD9;
        rom[241][21] = 16'h0016;
        rom[241][22] = 16'hFFCF;
        rom[241][23] = 16'h0004;
        rom[241][24] = 16'h0003;
        rom[241][25] = 16'hFFCE;
        rom[241][26] = 16'hFFFD;
        rom[241][27] = 16'h0004;
        rom[241][28] = 16'h000A;
        rom[241][29] = 16'hFFF2;
        rom[241][30] = 16'h0003;
        rom[241][31] = 16'h0003;
        rom[241][32] = 16'hFFEF;
        rom[241][33] = 16'hFFC3;
        rom[241][34] = 16'h000F;
        rom[241][35] = 16'hFFE4;
        rom[241][36] = 16'hFFDC;
        rom[241][37] = 16'h0000;
        rom[241][38] = 16'hFFF2;
        rom[241][39] = 16'hFFDA;
        rom[241][40] = 16'hFFFA;
        rom[241][41] = 16'hFFDC;
        rom[241][42] = 16'hFFF5;
        rom[241][43] = 16'h0037;
        rom[241][44] = 16'hFFF6;
        rom[241][45] = 16'h001C;
        rom[241][46] = 16'hFFB6;
        rom[241][47] = 16'hFFD5;
        rom[241][48] = 16'h0017;
        rom[241][49] = 16'h0002;
        rom[241][50] = 16'h001A;
        rom[241][51] = 16'hFFF5;
        rom[241][52] = 16'h0020;
        rom[241][53] = 16'h0008;
        rom[241][54] = 16'h001D;
        rom[241][55] = 16'hFFEA;
        rom[241][56] = 16'hFFF9;
        rom[241][57] = 16'hFFDB;
        rom[241][58] = 16'hFFD1;
        rom[241][59] = 16'h001A;
        rom[241][60] = 16'hFFF6;
        rom[241][61] = 16'hFFEE;
        rom[241][62] = 16'hFFEF;
        rom[241][63] = 16'hFFF5;
        rom[241][64] = 16'hFFE4;
        rom[241][65] = 16'hFFEA;
        rom[241][66] = 16'h000C;
        rom[241][67] = 16'h0024;
        rom[241][68] = 16'hFFD8;
        rom[241][69] = 16'h000D;
        rom[241][70] = 16'h0028;
        rom[241][71] = 16'h001A;
        rom[241][72] = 16'hFFEA;
        rom[241][73] = 16'h0007;
        rom[241][74] = 16'hFFCD;
        rom[241][75] = 16'h000B;
        rom[241][76] = 16'h0003;
        rom[241][77] = 16'hFFF4;
        rom[241][78] = 16'hFFEF;
        rom[241][79] = 16'hFFE1;
        rom[241][80] = 16'hFFE7;
        rom[241][81] = 16'h000F;
        rom[241][82] = 16'h0027;
        rom[241][83] = 16'h000C;
        rom[241][84] = 16'hFFC7;
        rom[241][85] = 16'h0002;
        rom[241][86] = 16'hFFEA;
        rom[241][87] = 16'hFFEA;
        rom[241][88] = 16'hFFEA;
        rom[241][89] = 16'h000A;
        rom[241][90] = 16'h0008;
        rom[241][91] = 16'hFFEA;
        rom[241][92] = 16'h0016;
        rom[241][93] = 16'hFFC4;
        rom[241][94] = 16'h0013;
        rom[241][95] = 16'hFFE1;
        rom[241][96] = 16'hFFDB;
        rom[241][97] = 16'hFFE8;
        rom[241][98] = 16'hFFFE;
        rom[241][99] = 16'hFFEB;
        rom[241][100] = 16'hFFF4;
        rom[241][101] = 16'h0008;
        rom[241][102] = 16'hFFF7;
        rom[241][103] = 16'hFFC4;
        rom[241][104] = 16'hFFF4;
        rom[241][105] = 16'hFF98;
        rom[241][106] = 16'h0007;
        rom[241][107] = 16'h0022;
        rom[241][108] = 16'hFFED;
        rom[241][109] = 16'hFFE4;
        rom[241][110] = 16'h000F;
        rom[241][111] = 16'hFFF5;
        rom[241][112] = 16'h001B;
        rom[241][113] = 16'hFFE5;
        rom[241][114] = 16'hFFD9;
        rom[241][115] = 16'hFFEC;
        rom[241][116] = 16'hFFDE;
        rom[241][117] = 16'h0011;
        rom[241][118] = 16'hFFDF;
        rom[241][119] = 16'h0002;
        rom[241][120] = 16'h000A;
        rom[241][121] = 16'hFFE7;
        rom[241][122] = 16'h0010;
        rom[241][123] = 16'h001B;
        rom[241][124] = 16'h0002;
        rom[241][125] = 16'h0003;
        rom[241][126] = 16'h0010;
        rom[241][127] = 16'h0006;
        rom[242][0] = 16'hFFEF;
        rom[242][1] = 16'h000F;
        rom[242][2] = 16'hFFEB;
        rom[242][3] = 16'h0006;
        rom[242][4] = 16'hFFD7;
        rom[242][5] = 16'hFFF4;
        rom[242][6] = 16'hFFF3;
        rom[242][7] = 16'h0021;
        rom[242][8] = 16'hFFC4;
        rom[242][9] = 16'hFFF6;
        rom[242][10] = 16'hFFFB;
        rom[242][11] = 16'hFFFE;
        rom[242][12] = 16'hFFC8;
        rom[242][13] = 16'h0024;
        rom[242][14] = 16'hFFFE;
        rom[242][15] = 16'hFFF4;
        rom[242][16] = 16'hFFFE;
        rom[242][17] = 16'h001F;
        rom[242][18] = 16'h000A;
        rom[242][19] = 16'hFFDF;
        rom[242][20] = 16'hFFED;
        rom[242][21] = 16'hFFB6;
        rom[242][22] = 16'hFFD2;
        rom[242][23] = 16'hFFF8;
        rom[242][24] = 16'hFFF7;
        rom[242][25] = 16'hFFCA;
        rom[242][26] = 16'hFFE3;
        rom[242][27] = 16'hFFBE;
        rom[242][28] = 16'hFFE5;
        rom[242][29] = 16'hFFFA;
        rom[242][30] = 16'hFFD2;
        rom[242][31] = 16'h0005;
        rom[242][32] = 16'hFFE5;
        rom[242][33] = 16'h001B;
        rom[242][34] = 16'hFFF9;
        rom[242][35] = 16'h0003;
        rom[242][36] = 16'hFFFB;
        rom[242][37] = 16'hFFC5;
        rom[242][38] = 16'hFFDF;
        rom[242][39] = 16'hFFF3;
        rom[242][40] = 16'h0016;
        rom[242][41] = 16'hFFB8;
        rom[242][42] = 16'hFFEA;
        rom[242][43] = 16'hFFEF;
        rom[242][44] = 16'hFFED;
        rom[242][45] = 16'hFFF8;
        rom[242][46] = 16'hFFEF;
        rom[242][47] = 16'h0022;
        rom[242][48] = 16'h0011;
        rom[242][49] = 16'h0011;
        rom[242][50] = 16'hFFEB;
        rom[242][51] = 16'hFFFE;
        rom[242][52] = 16'hFFFE;
        rom[242][53] = 16'h0017;
        rom[242][54] = 16'hFFFC;
        rom[242][55] = 16'hFFED;
        rom[242][56] = 16'h0002;
        rom[242][57] = 16'hFFE3;
        rom[242][58] = 16'h0017;
        rom[242][59] = 16'hFFE0;
        rom[242][60] = 16'hFFDF;
        rom[242][61] = 16'hFFF7;
        rom[242][62] = 16'h0008;
        rom[242][63] = 16'hFFF9;
        rom[242][64] = 16'hFFDF;
        rom[242][65] = 16'hFFEF;
        rom[242][66] = 16'hFFB5;
        rom[242][67] = 16'hFFD7;
        rom[242][68] = 16'hFFF7;
        rom[242][69] = 16'hFFCD;
        rom[242][70] = 16'hFFDB;
        rom[242][71] = 16'hFFED;
        rom[242][72] = 16'hFFDA;
        rom[242][73] = 16'hFFEF;
        rom[242][74] = 16'h0002;
        rom[242][75] = 16'hFFDC;
        rom[242][76] = 16'hFFE0;
        rom[242][77] = 16'h0005;
        rom[242][78] = 16'hFFAB;
        rom[242][79] = 16'hFFEF;
        rom[242][80] = 16'hFFFE;
        rom[242][81] = 16'h000F;
        rom[242][82] = 16'hFFFE;
        rom[242][83] = 16'hFFE8;
        rom[242][84] = 16'h000F;
        rom[242][85] = 16'hFFFC;
        rom[242][86] = 16'hFFFC;
        rom[242][87] = 16'h001B;
        rom[242][88] = 16'h002A;
        rom[242][89] = 16'h0019;
        rom[242][90] = 16'h0002;
        rom[242][91] = 16'hFFFE;
        rom[242][92] = 16'hFFFB;
        rom[242][93] = 16'hFFDF;
        rom[242][94] = 16'h0025;
        rom[242][95] = 16'hFFEF;
        rom[242][96] = 16'hFFE1;
        rom[242][97] = 16'h000C;
        rom[242][98] = 16'hFFF1;
        rom[242][99] = 16'hFFF9;
        rom[242][100] = 16'hFFB6;
        rom[242][101] = 16'hFFE3;
        rom[242][102] = 16'h0011;
        rom[242][103] = 16'hFFB5;
        rom[242][104] = 16'h001B;
        rom[242][105] = 16'h0010;
        rom[242][106] = 16'h0020;
        rom[242][107] = 16'hFFF3;
        rom[242][108] = 16'hFFC8;
        rom[242][109] = 16'hFFFC;
        rom[242][110] = 16'h000A;
        rom[242][111] = 16'hFFF4;
        rom[242][112] = 16'hFFD7;
        rom[242][113] = 16'hFFF9;
        rom[242][114] = 16'hFFE5;
        rom[242][115] = 16'hFFBA;
        rom[242][116] = 16'h0021;
        rom[242][117] = 16'hFFBE;
        rom[242][118] = 16'h000D;
        rom[242][119] = 16'hFFF9;
        rom[242][120] = 16'h0007;
        rom[242][121] = 16'hFFF7;
        rom[242][122] = 16'hFFD5;
        rom[242][123] = 16'h0014;
        rom[242][124] = 16'hFFF9;
        rom[242][125] = 16'hFFF4;
        rom[242][126] = 16'hFFF6;
        rom[242][127] = 16'hFFF4;
        rom[243][0] = 16'hFFDE;
        rom[243][1] = 16'hFFDE;
        rom[243][2] = 16'h0014;
        rom[243][3] = 16'hFFE7;
        rom[243][4] = 16'hFFFC;
        rom[243][5] = 16'h0016;
        rom[243][6] = 16'hFFFA;
        rom[243][7] = 16'hFFE6;
        rom[243][8] = 16'hFFE0;
        rom[243][9] = 16'h0004;
        rom[243][10] = 16'hFFE3;
        rom[243][11] = 16'h0013;
        rom[243][12] = 16'hFFF4;
        rom[243][13] = 16'h001C;
        rom[243][14] = 16'hFFF0;
        rom[243][15] = 16'h0016;
        rom[243][16] = 16'hFFFC;
        rom[243][17] = 16'h000D;
        rom[243][18] = 16'h0002;
        rom[243][19] = 16'h0004;
        rom[243][20] = 16'h001B;
        rom[243][21] = 16'hFFEF;
        rom[243][22] = 16'hFFBD;
        rom[243][23] = 16'hFFE2;
        rom[243][24] = 16'hFFEC;
        rom[243][25] = 16'h0002;
        rom[243][26] = 16'hFFE3;
        rom[243][27] = 16'h0014;
        rom[243][28] = 16'h0023;
        rom[243][29] = 16'h0028;
        rom[243][30] = 16'h000D;
        rom[243][31] = 16'hFFC6;
        rom[243][32] = 16'hFFED;
        rom[243][33] = 16'h0004;
        rom[243][34] = 16'h0007;
        rom[243][35] = 16'h0012;
        rom[243][36] = 16'hFFCB;
        rom[243][37] = 16'h000B;
        rom[243][38] = 16'hFFD4;
        rom[243][39] = 16'hFFDD;
        rom[243][40] = 16'h001B;
        rom[243][41] = 16'hFFFE;
        rom[243][42] = 16'hFFF5;
        rom[243][43] = 16'hFFF9;
        rom[243][44] = 16'hFFD8;
        rom[243][45] = 16'h0020;
        rom[243][46] = 16'hFFE6;
        rom[243][47] = 16'h000A;
        rom[243][48] = 16'hFFC6;
        rom[243][49] = 16'hFFDE;
        rom[243][50] = 16'hFFF0;
        rom[243][51] = 16'hFFCE;
        rom[243][52] = 16'h0018;
        rom[243][53] = 16'hFFED;
        rom[243][54] = 16'h002B;
        rom[243][55] = 16'h0016;
        rom[243][56] = 16'h0005;
        rom[243][57] = 16'hFFA8;
        rom[243][58] = 16'h0003;
        rom[243][59] = 16'h001B;
        rom[243][60] = 16'hFFFD;
        rom[243][61] = 16'h0027;
        rom[243][62] = 16'h0012;
        rom[243][63] = 16'hFFE3;
        rom[243][64] = 16'hFFFE;
        rom[243][65] = 16'hFFD2;
        rom[243][66] = 16'h0013;
        rom[243][67] = 16'hFFF9;
        rom[243][68] = 16'hFFE4;
        rom[243][69] = 16'hFFE0;
        rom[243][70] = 16'hFF9C;
        rom[243][71] = 16'hFFF2;
        rom[243][72] = 16'hFFFF;
        rom[243][73] = 16'hFFE1;
        rom[243][74] = 16'hFFBA;
        rom[243][75] = 16'hFFDC;
        rom[243][76] = 16'hFFFF;
        rom[243][77] = 16'h000D;
        rom[243][78] = 16'hFFF6;
        rom[243][79] = 16'hFFF4;
        rom[243][80] = 16'hFFE6;
        rom[243][81] = 16'h0018;
        rom[243][82] = 16'hFFD2;
        rom[243][83] = 16'hFFED;
        rom[243][84] = 16'hFFCC;
        rom[243][85] = 16'h0011;
        rom[243][86] = 16'h001C;
        rom[243][87] = 16'hFFFC;
        rom[243][88] = 16'hFFE4;
        rom[243][89] = 16'h001C;
        rom[243][90] = 16'hFFF6;
        rom[243][91] = 16'hFFEA;
        rom[243][92] = 16'hFFE7;
        rom[243][93] = 16'h001E;
        rom[243][94] = 16'h0020;
        rom[243][95] = 16'hFFE1;
        rom[243][96] = 16'hFFF7;
        rom[243][97] = 16'h0011;
        rom[243][98] = 16'h0001;
        rom[243][99] = 16'h001B;
        rom[243][100] = 16'hFFFD;
        rom[243][101] = 16'hFFFE;
        rom[243][102] = 16'hFFFF;
        rom[243][103] = 16'hFFC7;
        rom[243][104] = 16'hFFD7;
        rom[243][105] = 16'hFFF6;
        rom[243][106] = 16'h001D;
        rom[243][107] = 16'h0002;
        rom[243][108] = 16'h0045;
        rom[243][109] = 16'h000C;
        rom[243][110] = 16'h0027;
        rom[243][111] = 16'hFFFD;
        rom[243][112] = 16'h002F;
        rom[243][113] = 16'h0012;
        rom[243][114] = 16'h0003;
        rom[243][115] = 16'hFFE2;
        rom[243][116] = 16'hFFF9;
        rom[243][117] = 16'h001E;
        rom[243][118] = 16'h0009;
        rom[243][119] = 16'hFFDB;
        rom[243][120] = 16'h0014;
        rom[243][121] = 16'hFFFF;
        rom[243][122] = 16'h0007;
        rom[243][123] = 16'h0015;
        rom[243][124] = 16'h0014;
        rom[243][125] = 16'hFFE4;
        rom[243][126] = 16'h0016;
        rom[243][127] = 16'hFFF8;
        rom[244][0] = 16'hFFEC;
        rom[244][1] = 16'h0016;
        rom[244][2] = 16'h0004;
        rom[244][3] = 16'hFFFD;
        rom[244][4] = 16'h0051;
        rom[244][5] = 16'hFFEC;
        rom[244][6] = 16'hFFEF;
        rom[244][7] = 16'hFFE8;
        rom[244][8] = 16'h002C;
        rom[244][9] = 16'h0009;
        rom[244][10] = 16'hFFE7;
        rom[244][11] = 16'h001F;
        rom[244][12] = 16'h001E;
        rom[244][13] = 16'hFFF0;
        rom[244][14] = 16'h002B;
        rom[244][15] = 16'h0004;
        rom[244][16] = 16'hFFE7;
        rom[244][17] = 16'hFFEE;
        rom[244][18] = 16'hFFE1;
        rom[244][19] = 16'h0024;
        rom[244][20] = 16'h002F;
        rom[244][21] = 16'hFFF6;
        rom[244][22] = 16'h000C;
        rom[244][23] = 16'hFFEE;
        rom[244][24] = 16'h0011;
        rom[244][25] = 16'h000B;
        rom[244][26] = 16'hFFD2;
        rom[244][27] = 16'hFFEF;
        rom[244][28] = 16'hFFF6;
        rom[244][29] = 16'h002C;
        rom[244][30] = 16'h0007;
        rom[244][31] = 16'h0003;
        rom[244][32] = 16'hFFDC;
        rom[244][33] = 16'hFFCD;
        rom[244][34] = 16'h0011;
        rom[244][35] = 16'hFFF1;
        rom[244][36] = 16'hFFE3;
        rom[244][37] = 16'hFFEA;
        rom[244][38] = 16'h0028;
        rom[244][39] = 16'hFFCE;
        rom[244][40] = 16'h0035;
        rom[244][41] = 16'h0011;
        rom[244][42] = 16'hFFDF;
        rom[244][43] = 16'hFFE1;
        rom[244][44] = 16'hFFE0;
        rom[244][45] = 16'h0009;
        rom[244][46] = 16'hFFF9;
        rom[244][47] = 16'h0013;
        rom[244][48] = 16'hFFF9;
        rom[244][49] = 16'h001B;
        rom[244][50] = 16'h000D;
        rom[244][51] = 16'h0000;
        rom[244][52] = 16'h0008;
        rom[244][53] = 16'hFFFD;
        rom[244][54] = 16'h0000;
        rom[244][55] = 16'h0019;
        rom[244][56] = 16'h0022;
        rom[244][57] = 16'h001A;
        rom[244][58] = 16'h0009;
        rom[244][59] = 16'h000A;
        rom[244][60] = 16'hFFCD;
        rom[244][61] = 16'hFFF8;
        rom[244][62] = 16'h0023;
        rom[244][63] = 16'h000D;
        rom[244][64] = 16'hFFED;
        rom[244][65] = 16'h0003;
        rom[244][66] = 16'h0026;
        rom[244][67] = 16'h0023;
        rom[244][68] = 16'hFFE3;
        rom[244][69] = 16'h0037;
        rom[244][70] = 16'h002B;
        rom[244][71] = 16'hFFE7;
        rom[244][72] = 16'h0012;
        rom[244][73] = 16'h0011;
        rom[244][74] = 16'hFFF7;
        rom[244][75] = 16'hFFD4;
        rom[244][76] = 16'h0012;
        rom[244][77] = 16'hFFFF;
        rom[244][78] = 16'hFFDD;
        rom[244][79] = 16'h0024;
        rom[244][80] = 16'h0015;
        rom[244][81] = 16'hFFE3;
        rom[244][82] = 16'h0011;
        rom[244][83] = 16'h0037;
        rom[244][84] = 16'hFFEF;
        rom[244][85] = 16'h000F;
        rom[244][86] = 16'hFFF6;
        rom[244][87] = 16'h0010;
        rom[244][88] = 16'h000B;
        rom[244][89] = 16'h0002;
        rom[244][90] = 16'h0001;
        rom[244][91] = 16'hFFCD;
        rom[244][92] = 16'hFFCC;
        rom[244][93] = 16'hFFD2;
        rom[244][94] = 16'hFFCD;
        rom[244][95] = 16'hFFD5;
        rom[244][96] = 16'hFFE7;
        rom[244][97] = 16'hFFE5;
        rom[244][98] = 16'h0016;
        rom[244][99] = 16'hFFE6;
        rom[244][100] = 16'hFFDA;
        rom[244][101] = 16'hFFFE;
        rom[244][102] = 16'hFFF2;
        rom[244][103] = 16'h0016;
        rom[244][104] = 16'h0010;
        rom[244][105] = 16'h0015;
        rom[244][106] = 16'h002E;
        rom[244][107] = 16'h0011;
        rom[244][108] = 16'hFFB5;
        rom[244][109] = 16'hFFEF;
        rom[244][110] = 16'h0036;
        rom[244][111] = 16'hFFDB;
        rom[244][112] = 16'h000C;
        rom[244][113] = 16'hFFFE;
        rom[244][114] = 16'hFFD8;
        rom[244][115] = 16'hFFF4;
        rom[244][116] = 16'h0018;
        rom[244][117] = 16'h0000;
        rom[244][118] = 16'h000F;
        rom[244][119] = 16'h0012;
        rom[244][120] = 16'h002A;
        rom[244][121] = 16'hFFF7;
        rom[244][122] = 16'h002E;
        rom[244][123] = 16'hFFE6;
        rom[244][124] = 16'hFFF1;
        rom[244][125] = 16'h001F;
        rom[244][126] = 16'hFFFC;
        rom[244][127] = 16'hFFFD;
        rom[245][0] = 16'h000A;
        rom[245][1] = 16'h0012;
        rom[245][2] = 16'hFFFE;
        rom[245][3] = 16'hFFE6;
        rom[245][4] = 16'hFFD8;
        rom[245][5] = 16'hFFF3;
        rom[245][6] = 16'h002E;
        rom[245][7] = 16'hFFF4;
        rom[245][8] = 16'hFFEA;
        rom[245][9] = 16'hFFF0;
        rom[245][10] = 16'hFFFE;
        rom[245][11] = 16'h001A;
        rom[245][12] = 16'h002F;
        rom[245][13] = 16'h0019;
        rom[245][14] = 16'hFFF1;
        rom[245][15] = 16'hFFEE;
        rom[245][16] = 16'h000B;
        rom[245][17] = 16'h0019;
        rom[245][18] = 16'hFFB6;
        rom[245][19] = 16'h000C;
        rom[245][20] = 16'h000A;
        rom[245][21] = 16'hFFDA;
        rom[245][22] = 16'h0040;
        rom[245][23] = 16'h0017;
        rom[245][24] = 16'hFFE7;
        rom[245][25] = 16'h001F;
        rom[245][26] = 16'hFFDF;
        rom[245][27] = 16'h001E;
        rom[245][28] = 16'h000C;
        rom[245][29] = 16'h0010;
        rom[245][30] = 16'hFFE0;
        rom[245][31] = 16'h0028;
        rom[245][32] = 16'hFFF5;
        rom[245][33] = 16'h0002;
        rom[245][34] = 16'h001E;
        rom[245][35] = 16'h0026;
        rom[245][36] = 16'h0013;
        rom[245][37] = 16'hFFD7;
        rom[245][38] = 16'hFFE3;
        rom[245][39] = 16'h0002;
        rom[245][40] = 16'h000D;
        rom[245][41] = 16'hFFFE;
        rom[245][42] = 16'h0011;
        rom[245][43] = 16'h0020;
        rom[245][44] = 16'h0017;
        rom[245][45] = 16'h0026;
        rom[245][46] = 16'hFFF9;
        rom[245][47] = 16'h0011;
        rom[245][48] = 16'hFFF8;
        rom[245][49] = 16'hFFE3;
        rom[245][50] = 16'h0005;
        rom[245][51] = 16'hFFF0;
        rom[245][52] = 16'h001E;
        rom[245][53] = 16'hFFBC;
        rom[245][54] = 16'hFFC7;
        rom[245][55] = 16'h001A;
        rom[245][56] = 16'hFFE9;
        rom[245][57] = 16'h0009;
        rom[245][58] = 16'hFFF4;
        rom[245][59] = 16'hFFFC;
        rom[245][60] = 16'h0003;
        rom[245][61] = 16'h0003;
        rom[245][62] = 16'h0002;
        rom[245][63] = 16'hFFF5;
        rom[245][64] = 16'hFFF4;
        rom[245][65] = 16'hFFE4;
        rom[245][66] = 16'hFFE1;
        rom[245][67] = 16'hFFDC;
        rom[245][68] = 16'hFFB0;
        rom[245][69] = 16'hFFF5;
        rom[245][70] = 16'hFFBA;
        rom[245][71] = 16'h0015;
        rom[245][72] = 16'hFFD7;
        rom[245][73] = 16'hFFCF;
        rom[245][74] = 16'hFFCC;
        rom[245][75] = 16'hFFCE;
        rom[245][76] = 16'hFFF7;
        rom[245][77] = 16'hFFEA;
        rom[245][78] = 16'hFFE2;
        rom[245][79] = 16'h000A;
        rom[245][80] = 16'h0017;
        rom[245][81] = 16'h001F;
        rom[245][82] = 16'hFFF3;
        rom[245][83] = 16'h001E;
        rom[245][84] = 16'h000F;
        rom[245][85] = 16'hFFDE;
        rom[245][86] = 16'hFFCA;
        rom[245][87] = 16'h000C;
        rom[245][88] = 16'hFFF0;
        rom[245][89] = 16'hFFB4;
        rom[245][90] = 16'hFFF9;
        rom[245][91] = 16'hFFF2;
        rom[245][92] = 16'hFFE0;
        rom[245][93] = 16'hFFE9;
        rom[245][94] = 16'hFFFD;
        rom[245][95] = 16'h0003;
        rom[245][96] = 16'hFFF4;
        rom[245][97] = 16'hFFDF;
        rom[245][98] = 16'hFFFC;
        rom[245][99] = 16'h000B;
        rom[245][100] = 16'hFFF4;
        rom[245][101] = 16'h001A;
        rom[245][102] = 16'h002D;
        rom[245][103] = 16'h0038;
        rom[245][104] = 16'h0015;
        rom[245][105] = 16'h000C;
        rom[245][106] = 16'h0002;
        rom[245][107] = 16'hFFE6;
        rom[245][108] = 16'h0014;
        rom[245][109] = 16'hFFF0;
        rom[245][110] = 16'h0016;
        rom[245][111] = 16'h0012;
        rom[245][112] = 16'h0016;
        rom[245][113] = 16'h0011;
        rom[245][114] = 16'h0029;
        rom[245][115] = 16'h0000;
        rom[245][116] = 16'h0045;
        rom[245][117] = 16'hFFD7;
        rom[245][118] = 16'hFFF1;
        rom[245][119] = 16'h0007;
        rom[245][120] = 16'hFFDB;
        rom[245][121] = 16'hFFEA;
        rom[245][122] = 16'hFFCA;
        rom[245][123] = 16'hFFEE;
        rom[245][124] = 16'hFFBE;
        rom[245][125] = 16'hFFB5;
        rom[245][126] = 16'h000B;
        rom[245][127] = 16'hFFF9;
        rom[246][0] = 16'hFFF4;
        rom[246][1] = 16'hFFCE;
        rom[246][2] = 16'hFFF7;
        rom[246][3] = 16'hFFFE;
        rom[246][4] = 16'hFFF3;
        rom[246][5] = 16'h0005;
        rom[246][6] = 16'hFFF9;
        rom[246][7] = 16'hFFBB;
        rom[246][8] = 16'hFFBD;
        rom[246][9] = 16'hFFD5;
        rom[246][10] = 16'h0006;
        rom[246][11] = 16'hFFE8;
        rom[246][12] = 16'h0000;
        rom[246][13] = 16'hFFEA;
        rom[246][14] = 16'hFFEE;
        rom[246][15] = 16'hFFEC;
        rom[246][16] = 16'h0014;
        rom[246][17] = 16'hFFC5;
        rom[246][18] = 16'h0002;
        rom[246][19] = 16'h001F;
        rom[246][20] = 16'h0007;
        rom[246][21] = 16'hFFDF;
        rom[246][22] = 16'hFFEF;
        rom[246][23] = 16'hFFC3;
        rom[246][24] = 16'hFFC3;
        rom[246][25] = 16'hFFEB;
        rom[246][26] = 16'h0015;
        rom[246][27] = 16'h000C;
        rom[246][28] = 16'h0007;
        rom[246][29] = 16'hFFC9;
        rom[246][30] = 16'hFFE8;
        rom[246][31] = 16'hFFB5;
        rom[246][32] = 16'h0011;
        rom[246][33] = 16'hFFC4;
        rom[246][34] = 16'hFFD6;
        rom[246][35] = 16'hFFE4;
        rom[246][36] = 16'hFFE9;
        rom[246][37] = 16'hFFE7;
        rom[246][38] = 16'hFF98;
        rom[246][39] = 16'h001A;
        rom[246][40] = 16'hFFE1;
        rom[246][41] = 16'h0007;
        rom[246][42] = 16'hFFFC;
        rom[246][43] = 16'hFFF9;
        rom[246][44] = 16'h0012;
        rom[246][45] = 16'h0015;
        rom[246][46] = 16'h0038;
        rom[246][47] = 16'hFFCD;
        rom[246][48] = 16'hFFF7;
        rom[246][49] = 16'h0028;
        rom[246][50] = 16'h0011;
        rom[246][51] = 16'h0015;
        rom[246][52] = 16'h000D;
        rom[246][53] = 16'h000C;
        rom[246][54] = 16'h0002;
        rom[246][55] = 16'hFFC3;
        rom[246][56] = 16'h0009;
        rom[246][57] = 16'hFFD2;
        rom[246][58] = 16'hFFBB;
        rom[246][59] = 16'hFFF3;
        rom[246][60] = 16'h0029;
        rom[246][61] = 16'hFFF9;
        rom[246][62] = 16'h0018;
        rom[246][63] = 16'hFFF2;
        rom[246][64] = 16'hFFCC;
        rom[246][65] = 16'hFFDC;
        rom[246][66] = 16'hFFE9;
        rom[246][67] = 16'h0000;
        rom[246][68] = 16'h000F;
        rom[246][69] = 16'h000C;
        rom[246][70] = 16'hFFB0;
        rom[246][71] = 16'h0006;
        rom[246][72] = 16'h0011;
        rom[246][73] = 16'hFFDC;
        rom[246][74] = 16'hFFE1;
        rom[246][75] = 16'hFFE5;
        rom[246][76] = 16'hFFC4;
        rom[246][77] = 16'hFFF9;
        rom[246][78] = 16'hFFF4;
        rom[246][79] = 16'hFFC2;
        rom[246][80] = 16'hFFE6;
        rom[246][81] = 16'h0012;
        rom[246][82] = 16'hFFD6;
        rom[246][83] = 16'hFFBF;
        rom[246][84] = 16'h0007;
        rom[246][85] = 16'h000D;
        rom[246][86] = 16'h001F;
        rom[246][87] = 16'h001B;
        rom[246][88] = 16'hFFEA;
        rom[246][89] = 16'h0019;
        rom[246][90] = 16'h0004;
        rom[246][91] = 16'h0009;
        rom[246][92] = 16'hFFD0;
        rom[246][93] = 16'h000B;
        rom[246][94] = 16'hFFE1;
        rom[246][95] = 16'hFFFF;
        rom[246][96] = 16'h0011;
        rom[246][97] = 16'h0019;
        rom[246][98] = 16'h001F;
        rom[246][99] = 16'h003E;
        rom[246][100] = 16'h000F;
        rom[246][101] = 16'h0002;
        rom[246][102] = 16'h0001;
        rom[246][103] = 16'hFFF0;
        rom[246][104] = 16'hFFF6;
        rom[246][105] = 16'h0024;
        rom[246][106] = 16'hFFD2;
        rom[246][107] = 16'h0006;
        rom[246][108] = 16'h0046;
        rom[246][109] = 16'h001C;
        rom[246][110] = 16'hFFEE;
        rom[246][111] = 16'h001B;
        rom[246][112] = 16'h0019;
        rom[246][113] = 16'hFFEC;
        rom[246][114] = 16'h000D;
        rom[246][115] = 16'hFFC3;
        rom[246][116] = 16'hFFAF;
        rom[246][117] = 16'h0024;
        rom[246][118] = 16'h0013;
        rom[246][119] = 16'hFFF7;
        rom[246][120] = 16'h0002;
        rom[246][121] = 16'h001C;
        rom[246][122] = 16'hFFFA;
        rom[246][123] = 16'h0002;
        rom[246][124] = 16'h000C;
        rom[246][125] = 16'h0000;
        rom[246][126] = 16'h0008;
        rom[246][127] = 16'h0011;
        rom[247][0] = 16'h0024;
        rom[247][1] = 16'hFFEA;
        rom[247][2] = 16'hFF9B;
        rom[247][3] = 16'h000A;
        rom[247][4] = 16'hFFFB;
        rom[247][5] = 16'h0016;
        rom[247][6] = 16'hFFE9;
        rom[247][7] = 16'h0002;
        rom[247][8] = 16'h0009;
        rom[247][9] = 16'hFFEA;
        rom[247][10] = 16'h0015;
        rom[247][11] = 16'hFFCD;
        rom[247][12] = 16'h0015;
        rom[247][13] = 16'h000C;
        rom[247][14] = 16'hFFF3;
        rom[247][15] = 16'h0009;
        rom[247][16] = 16'hFFF9;
        rom[247][17] = 16'h0012;
        rom[247][18] = 16'hFFEB;
        rom[247][19] = 16'h0018;
        rom[247][20] = 16'hFFDA;
        rom[247][21] = 16'h001E;
        rom[247][22] = 16'h000B;
        rom[247][23] = 16'h004B;
        rom[247][24] = 16'hFFA2;
        rom[247][25] = 16'hFFB0;
        rom[247][26] = 16'h0006;
        rom[247][27] = 16'hFFE3;
        rom[247][28] = 16'hFFF4;
        rom[247][29] = 16'hFFE1;
        rom[247][30] = 16'h0029;
        rom[247][31] = 16'h0004;
        rom[247][32] = 16'hFFEC;
        rom[247][33] = 16'h002A;
        rom[247][34] = 16'h0000;
        rom[247][35] = 16'h0007;
        rom[247][36] = 16'hFFDB;
        rom[247][37] = 16'hFFCE;
        rom[247][38] = 16'h0011;
        rom[247][39] = 16'h0029;
        rom[247][40] = 16'hFFFF;
        rom[247][41] = 16'h0024;
        rom[247][42] = 16'h000B;
        rom[247][43] = 16'hFFEA;
        rom[247][44] = 16'h0026;
        rom[247][45] = 16'h001A;
        rom[247][46] = 16'h0004;
        rom[247][47] = 16'h001C;
        rom[247][48] = 16'h0002;
        rom[247][49] = 16'hFFD2;
        rom[247][50] = 16'hFFFB;
        rom[247][51] = 16'h000A;
        rom[247][52] = 16'h0020;
        rom[247][53] = 16'h0006;
        rom[247][54] = 16'h000F;
        rom[247][55] = 16'hFFF7;
        rom[247][56] = 16'h000D;
        rom[247][57] = 16'h0036;
        rom[247][58] = 16'hFFF9;
        rom[247][59] = 16'hFFBC;
        rom[247][60] = 16'h0006;
        rom[247][61] = 16'hFFEE;
        rom[247][62] = 16'hFFEF;
        rom[247][63] = 16'hFFE2;
        rom[247][64] = 16'hFFC8;
        rom[247][65] = 16'hFFD9;
        rom[247][66] = 16'hFFF1;
        rom[247][67] = 16'hFFFE;
        rom[247][68] = 16'hFFEE;
        rom[247][69] = 16'hFFF9;
        rom[247][70] = 16'hFFFB;
        rom[247][71] = 16'hFFF5;
        rom[247][72] = 16'h0017;
        rom[247][73] = 16'h0003;
        rom[247][74] = 16'h001B;
        rom[247][75] = 16'hFFC8;
        rom[247][76] = 16'hFF9D;
        rom[247][77] = 16'h001F;
        rom[247][78] = 16'h003D;
        rom[247][79] = 16'h001C;
        rom[247][80] = 16'hFFF9;
        rom[247][81] = 16'h000C;
        rom[247][82] = 16'h0003;
        rom[247][83] = 16'h002A;
        rom[247][84] = 16'hFFF3;
        rom[247][85] = 16'h0024;
        rom[247][86] = 16'hFFE3;
        rom[247][87] = 16'h0014;
        rom[247][88] = 16'hFFFE;
        rom[247][89] = 16'h0035;
        rom[247][90] = 16'hFFF3;
        rom[247][91] = 16'hFFF2;
        rom[247][92] = 16'hFF99;
        rom[247][93] = 16'h0027;
        rom[247][94] = 16'h0009;
        rom[247][95] = 16'h0011;
        rom[247][96] = 16'h0010;
        rom[247][97] = 16'h000A;
        rom[247][98] = 16'h000D;
        rom[247][99] = 16'h0003;
        rom[247][100] = 16'hFFF0;
        rom[247][101] = 16'hFFEE;
        rom[247][102] = 16'hFF9D;
        rom[247][103] = 16'hFFE1;
        rom[247][104] = 16'h0002;
        rom[247][105] = 16'h0011;
        rom[247][106] = 16'hFFC1;
        rom[247][107] = 16'h0027;
        rom[247][108] = 16'hFFE4;
        rom[247][109] = 16'h0011;
        rom[247][110] = 16'hFFF5;
        rom[247][111] = 16'h0012;
        rom[247][112] = 16'hFFF4;
        rom[247][113] = 16'h0021;
        rom[247][114] = 16'hFFF1;
        rom[247][115] = 16'hFFF4;
        rom[247][116] = 16'h0032;
        rom[247][117] = 16'h0007;
        rom[247][118] = 16'h0017;
        rom[247][119] = 16'h001E;
        rom[247][120] = 16'h002D;
        rom[247][121] = 16'h001A;
        rom[247][122] = 16'hFFF0;
        rom[247][123] = 16'hFFEC;
        rom[247][124] = 16'h0029;
        rom[247][125] = 16'h0032;
        rom[247][126] = 16'h0002;
        rom[247][127] = 16'h000F;
        rom[248][0] = 16'hFFF5;
        rom[248][1] = 16'hFFD3;
        rom[248][2] = 16'hFFFF;
        rom[248][3] = 16'hFFCD;
        rom[248][4] = 16'hFFCC;
        rom[248][5] = 16'h0000;
        rom[248][6] = 16'h0003;
        rom[248][7] = 16'h0005;
        rom[248][8] = 16'h000D;
        rom[248][9] = 16'hFFBA;
        rom[248][10] = 16'h001C;
        rom[248][11] = 16'h000C;
        rom[248][12] = 16'hFFF6;
        rom[248][13] = 16'h0012;
        rom[248][14] = 16'hFFCD;
        rom[248][15] = 16'h0022;
        rom[248][16] = 16'h000A;
        rom[248][17] = 16'h0024;
        rom[248][18] = 16'hFFC0;
        rom[248][19] = 16'hFFE6;
        rom[248][20] = 16'hFFCD;
        rom[248][21] = 16'h0009;
        rom[248][22] = 16'hFFF1;
        rom[248][23] = 16'hFFE4;
        rom[248][24] = 16'hFFDC;
        rom[248][25] = 16'hFFF9;
        rom[248][26] = 16'hFFD5;
        rom[248][27] = 16'h000C;
        rom[248][28] = 16'h0048;
        rom[248][29] = 16'h0001;
        rom[248][30] = 16'hFFF7;
        rom[248][31] = 16'h0027;
        rom[248][32] = 16'hFFEA;
        rom[248][33] = 16'hFFFF;
        rom[248][34] = 16'hFFF3;
        rom[248][35] = 16'h0012;
        rom[248][36] = 16'hFFE4;
        rom[248][37] = 16'hFFC1;
        rom[248][38] = 16'hFFEC;
        rom[248][39] = 16'hFFCE;
        rom[248][40] = 16'h000C;
        rom[248][41] = 16'hFFDD;
        rom[248][42] = 16'h0007;
        rom[248][43] = 16'h002A;
        rom[248][44] = 16'hFFF1;
        rom[248][45] = 16'h0016;
        rom[248][46] = 16'hFFBE;
        rom[248][47] = 16'h000B;
        rom[248][48] = 16'hFFE5;
        rom[248][49] = 16'hFFE4;
        rom[248][50] = 16'h0000;
        rom[248][51] = 16'hFFE5;
        rom[248][52] = 16'h0016;
        rom[248][53] = 16'h000E;
        rom[248][54] = 16'hFFFE;
        rom[248][55] = 16'hFFE5;
        rom[248][56] = 16'h0013;
        rom[248][57] = 16'hFFEA;
        rom[248][58] = 16'hFFFE;
        rom[248][59] = 16'hFFE6;
        rom[248][60] = 16'hFFDC;
        rom[248][61] = 16'h0018;
        rom[248][62] = 16'hFFF9;
        rom[248][63] = 16'hFFEE;
        rom[248][64] = 16'h000D;
        rom[248][65] = 16'h0009;
        rom[248][66] = 16'hFFEA;
        rom[248][67] = 16'h0008;
        rom[248][68] = 16'hFFFA;
        rom[248][69] = 16'h0011;
        rom[248][70] = 16'hFFF1;
        rom[248][71] = 16'h0011;
        rom[248][72] = 16'hFFEB;
        rom[248][73] = 16'hFFF8;
        rom[248][74] = 16'h0032;
        rom[248][75] = 16'h0004;
        rom[248][76] = 16'h001C;
        rom[248][77] = 16'h000A;
        rom[248][78] = 16'hFFCA;
        rom[248][79] = 16'hFFEA;
        rom[248][80] = 16'h0006;
        rom[248][81] = 16'hFFF8;
        rom[248][82] = 16'h0006;
        rom[248][83] = 16'hFFEC;
        rom[248][84] = 16'hFFD7;
        rom[248][85] = 16'h0019;
        rom[248][86] = 16'hFFEF;
        rom[248][87] = 16'h000C;
        rom[248][88] = 16'hFFBC;
        rom[248][89] = 16'h001B;
        rom[248][90] = 16'hFFF8;
        rom[248][91] = 16'h0018;
        rom[248][92] = 16'h0016;
        rom[248][93] = 16'hFFF7;
        rom[248][94] = 16'h0046;
        rom[248][95] = 16'hFFDD;
        rom[248][96] = 16'hFFE9;
        rom[248][97] = 16'hFFE8;
        rom[248][98] = 16'h000D;
        rom[248][99] = 16'h001A;
        rom[248][100] = 16'h002A;
        rom[248][101] = 16'hFFD4;
        rom[248][102] = 16'h001E;
        rom[248][103] = 16'h000C;
        rom[248][104] = 16'hFFFA;
        rom[248][105] = 16'hFFD0;
        rom[248][106] = 16'h003D;
        rom[248][107] = 16'h0011;
        rom[248][108] = 16'h0032;
        rom[248][109] = 16'hFFED;
        rom[248][110] = 16'h001B;
        rom[248][111] = 16'h0018;
        rom[248][112] = 16'h0001;
        rom[248][113] = 16'hFFE2;
        rom[248][114] = 16'h0014;
        rom[248][115] = 16'hFFE1;
        rom[248][116] = 16'hFFFA;
        rom[248][117] = 16'hFFCD;
        rom[248][118] = 16'hFFE3;
        rom[248][119] = 16'hFFDC;
        rom[248][120] = 16'h0019;
        rom[248][121] = 16'h0006;
        rom[248][122] = 16'h000A;
        rom[248][123] = 16'h000C;
        rom[248][124] = 16'hFFF6;
        rom[248][125] = 16'hFFFE;
        rom[248][126] = 16'h001F;
        rom[248][127] = 16'h0016;
        rom[249][0] = 16'hFFE1;
        rom[249][1] = 16'h001A;
        rom[249][2] = 16'h0008;
        rom[249][3] = 16'hFFDD;
        rom[249][4] = 16'hFFDC;
        rom[249][5] = 16'h000E;
        rom[249][6] = 16'h001B;
        rom[249][7] = 16'hFFC8;
        rom[249][8] = 16'hFFF9;
        rom[249][9] = 16'hFFBA;
        rom[249][10] = 16'hFFF0;
        rom[249][11] = 16'hFFF2;
        rom[249][12] = 16'h001D;
        rom[249][13] = 16'hFFD8;
        rom[249][14] = 16'hFFF9;
        rom[249][15] = 16'h0032;
        rom[249][16] = 16'h0001;
        rom[249][17] = 16'hFFCD;
        rom[249][18] = 16'h0008;
        rom[249][19] = 16'h0028;
        rom[249][20] = 16'hFFFE;
        rom[249][21] = 16'hFFE7;
        rom[249][22] = 16'hFFF1;
        rom[249][23] = 16'hFFF7;
        rom[249][24] = 16'hFFD8;
        rom[249][25] = 16'h001A;
        rom[249][26] = 16'h0004;
        rom[249][27] = 16'hFFFF;
        rom[249][28] = 16'h0014;
        rom[249][29] = 16'h0016;
        rom[249][30] = 16'hFFD2;
        rom[249][31] = 16'hFFB2;
        rom[249][32] = 16'hFFFD;
        rom[249][33] = 16'hFFC8;
        rom[249][34] = 16'hFFD9;
        rom[249][35] = 16'h0012;
        rom[249][36] = 16'hFFFA;
        rom[249][37] = 16'h001A;
        rom[249][38] = 16'hFFB4;
        rom[249][39] = 16'h001A;
        rom[249][40] = 16'hFFA9;
        rom[249][41] = 16'h0012;
        rom[249][42] = 16'hFFFE;
        rom[249][43] = 16'h001B;
        rom[249][44] = 16'hFFF8;
        rom[249][45] = 16'h0034;
        rom[249][46] = 16'h0002;
        rom[249][47] = 16'h0009;
        rom[249][48] = 16'hFFF6;
        rom[249][49] = 16'h0018;
        rom[249][50] = 16'hFFD4;
        rom[249][51] = 16'hFFCC;
        rom[249][52] = 16'h0000;
        rom[249][53] = 16'hFFEB;
        rom[249][54] = 16'h0000;
        rom[249][55] = 16'hFFDF;
        rom[249][56] = 16'hFFFB;
        rom[249][57] = 16'hFFC3;
        rom[249][58] = 16'hFFED;
        rom[249][59] = 16'h0021;
        rom[249][60] = 16'h0010;
        rom[249][61] = 16'h0006;
        rom[249][62] = 16'h0034;
        rom[249][63] = 16'hFFE7;
        rom[249][64] = 16'hFFF8;
        rom[249][65] = 16'hFFF4;
        rom[249][66] = 16'hFFF8;
        rom[249][67] = 16'h0012;
        rom[249][68] = 16'hFFED;
        rom[249][69] = 16'hFFF9;
        rom[249][70] = 16'hFFEF;
        rom[249][71] = 16'h000D;
        rom[249][72] = 16'hFFD8;
        rom[249][73] = 16'h0001;
        rom[249][74] = 16'hFFB4;
        rom[249][75] = 16'hFFBB;
        rom[249][76] = 16'hFFFE;
        rom[249][77] = 16'hFFBB;
        rom[249][78] = 16'hFFEC;
        rom[249][79] = 16'hFFF0;
        rom[249][80] = 16'h0007;
        rom[249][81] = 16'h0036;
        rom[249][82] = 16'h0017;
        rom[249][83] = 16'hFFDC;
        rom[249][84] = 16'h000B;
        rom[249][85] = 16'hFFB1;
        rom[249][86] = 16'h0011;
        rom[249][87] = 16'hFFC5;
        rom[249][88] = 16'hFFF5;
        rom[249][89] = 16'h0025;
        rom[249][90] = 16'hFFFB;
        rom[249][91] = 16'h0016;
        rom[249][92] = 16'hFFC4;
        rom[249][93] = 16'h000C;
        rom[249][94] = 16'hFFCE;
        rom[249][95] = 16'h0009;
        rom[249][96] = 16'h0002;
        rom[249][97] = 16'h0019;
        rom[249][98] = 16'h000F;
        rom[249][99] = 16'h0040;
        rom[249][100] = 16'h0007;
        rom[249][101] = 16'hFFF0;
        rom[249][102] = 16'h0014;
        rom[249][103] = 16'hFFCF;
        rom[249][104] = 16'hFFDC;
        rom[249][105] = 16'h000E;
        rom[249][106] = 16'h000E;
        rom[249][107] = 16'h001C;
        rom[249][108] = 16'h0004;
        rom[249][109] = 16'h000D;
        rom[249][110] = 16'h0017;
        rom[249][111] = 16'h0029;
        rom[249][112] = 16'h0005;
        rom[249][113] = 16'h0004;
        rom[249][114] = 16'hFFFE;
        rom[249][115] = 16'hFFD0;
        rom[249][116] = 16'hFFFD;
        rom[249][117] = 16'h0039;
        rom[249][118] = 16'hFFFF;
        rom[249][119] = 16'h001B;
        rom[249][120] = 16'hFFE5;
        rom[249][121] = 16'hFFE6;
        rom[249][122] = 16'hFFEA;
        rom[249][123] = 16'hFFC2;
        rom[249][124] = 16'h001B;
        rom[249][125] = 16'hFFE6;
        rom[249][126] = 16'hFFD7;
        rom[249][127] = 16'h0003;
        rom[250][0] = 16'h0000;
        rom[250][1] = 16'h0013;
        rom[250][2] = 16'hFFFE;
        rom[250][3] = 16'hFFD3;
        rom[250][4] = 16'h0022;
        rom[250][5] = 16'h001F;
        rom[250][6] = 16'hFFFB;
        rom[250][7] = 16'h0023;
        rom[250][8] = 16'h001A;
        rom[250][9] = 16'h0004;
        rom[250][10] = 16'hFFD2;
        rom[250][11] = 16'h0019;
        rom[250][12] = 16'hFFF4;
        rom[250][13] = 16'hFFB5;
        rom[250][14] = 16'h0002;
        rom[250][15] = 16'h0013;
        rom[250][16] = 16'h0003;
        rom[250][17] = 16'hFFDE;
        rom[250][18] = 16'h001F;
        rom[250][19] = 16'h0010;
        rom[250][20] = 16'hFFDE;
        rom[250][21] = 16'hFFFA;
        rom[250][22] = 16'h0001;
        rom[250][23] = 16'h0000;
        rom[250][24] = 16'h0003;
        rom[250][25] = 16'hFFF9;
        rom[250][26] = 16'hFFF6;
        rom[250][27] = 16'hFFC5;
        rom[250][28] = 16'hFFE8;
        rom[250][29] = 16'hFFE1;
        rom[250][30] = 16'hFFEF;
        rom[250][31] = 16'hFFF4;
        rom[250][32] = 16'h000E;
        rom[250][33] = 16'h000F;
        rom[250][34] = 16'h000B;
        rom[250][35] = 16'hFFC3;
        rom[250][36] = 16'h0019;
        rom[250][37] = 16'hFFC4;
        rom[250][38] = 16'h0016;
        rom[250][39] = 16'hFFDB;
        rom[250][40] = 16'hFFC8;
        rom[250][41] = 16'h0012;
        rom[250][42] = 16'hFFEC;
        rom[250][43] = 16'h000C;
        rom[250][44] = 16'hFFD5;
        rom[250][45] = 16'hFFC8;
        rom[250][46] = 16'h0003;
        rom[250][47] = 16'h0010;
        rom[250][48] = 16'h0014;
        rom[250][49] = 16'h001D;
        rom[250][50] = 16'h000A;
        rom[250][51] = 16'hFFD5;
        rom[250][52] = 16'h002B;
        rom[250][53] = 16'hFFE4;
        rom[250][54] = 16'hFFBF;
        rom[250][55] = 16'h0016;
        rom[250][56] = 16'hFFD7;
        rom[250][57] = 16'hFFE7;
        rom[250][58] = 16'h0016;
        rom[250][59] = 16'hFFE1;
        rom[250][60] = 16'hFFEC;
        rom[250][61] = 16'hFFE6;
        rom[250][62] = 16'hFFEA;
        rom[250][63] = 16'h0007;
        rom[250][64] = 16'h002F;
        rom[250][65] = 16'hFFF8;
        rom[250][66] = 16'h002F;
        rom[250][67] = 16'h0024;
        rom[250][68] = 16'hFFF6;
        rom[250][69] = 16'hFFF4;
        rom[250][70] = 16'h0016;
        rom[250][71] = 16'h0019;
        rom[250][72] = 16'hFFD3;
        rom[250][73] = 16'hFFEA;
        rom[250][74] = 16'hFFCC;
        rom[250][75] = 16'h0033;
        rom[250][76] = 16'h001B;
        rom[250][77] = 16'hFFE3;
        rom[250][78] = 16'hFFEA;
        rom[250][79] = 16'h0022;
        rom[250][80] = 16'h0004;
        rom[250][81] = 16'h001C;
        rom[250][82] = 16'h0019;
        rom[250][83] = 16'hFFD8;
        rom[250][84] = 16'h0012;
        rom[250][85] = 16'h001B;
        rom[250][86] = 16'hFFD4;
        rom[250][87] = 16'h0027;
        rom[250][88] = 16'hFFE5;
        rom[250][89] = 16'hFFC3;
        rom[250][90] = 16'h0017;
        rom[250][91] = 16'h001B;
        rom[250][92] = 16'hFFF3;
        rom[250][93] = 16'hFFE7;
        rom[250][94] = 16'hFFE0;
        rom[250][95] = 16'h0002;
        rom[250][96] = 16'h0019;
        rom[250][97] = 16'h0008;
        rom[250][98] = 16'hFFE5;
        rom[250][99] = 16'h0018;
        rom[250][100] = 16'hFFDE;
        rom[250][101] = 16'h0008;
        rom[250][102] = 16'hFFF4;
        rom[250][103] = 16'h001E;
        rom[250][104] = 16'h000C;
        rom[250][105] = 16'h000D;
        rom[250][106] = 16'h000A;
        rom[250][107] = 16'h0015;
        rom[250][108] = 16'hFFFA;
        rom[250][109] = 16'hFFEF;
        rom[250][110] = 16'h0032;
        rom[250][111] = 16'h0018;
        rom[250][112] = 16'hFFE8;
        rom[250][113] = 16'hFFF0;
        rom[250][114] = 16'h0002;
        rom[250][115] = 16'hFFE3;
        rom[250][116] = 16'h003E;
        rom[250][117] = 16'h0020;
        rom[250][118] = 16'hFFF7;
        rom[250][119] = 16'hFFF6;
        rom[250][120] = 16'hFFF2;
        rom[250][121] = 16'hFFEC;
        rom[250][122] = 16'h000F;
        rom[250][123] = 16'h000F;
        rom[250][124] = 16'hFFF4;
        rom[250][125] = 16'h0002;
        rom[250][126] = 16'hFFF6;
        rom[250][127] = 16'h0029;
        rom[251][0] = 16'h0024;
        rom[251][1] = 16'hFFEA;
        rom[251][2] = 16'h000A;
        rom[251][3] = 16'hFFEA;
        rom[251][4] = 16'hFFE2;
        rom[251][5] = 16'hFFFB;
        rom[251][6] = 16'hFFD1;
        rom[251][7] = 16'hFFDA;
        rom[251][8] = 16'h000E;
        rom[251][9] = 16'h001F;
        rom[251][10] = 16'hFFD3;
        rom[251][11] = 16'h0026;
        rom[251][12] = 16'h002E;
        rom[251][13] = 16'h0000;
        rom[251][14] = 16'hFFF1;
        rom[251][15] = 16'hFFFE;
        rom[251][16] = 16'hFFE3;
        rom[251][17] = 16'h0005;
        rom[251][18] = 16'hFFF4;
        rom[251][19] = 16'h0016;
        rom[251][20] = 16'h000C;
        rom[251][21] = 16'h000F;
        rom[251][22] = 16'h002F;
        rom[251][23] = 16'hFFD5;
        rom[251][24] = 16'hFFDC;
        rom[251][25] = 16'hFFEA;
        rom[251][26] = 16'hFFC6;
        rom[251][27] = 16'hFFF7;
        rom[251][28] = 16'h001F;
        rom[251][29] = 16'h001A;
        rom[251][30] = 16'hFFE3;
        rom[251][31] = 16'hFFEB;
        rom[251][32] = 16'h001E;
        rom[251][33] = 16'hFFF2;
        rom[251][34] = 16'hFFC8;
        rom[251][35] = 16'hFFFB;
        rom[251][36] = 16'hFFEA;
        rom[251][37] = 16'hFFEF;
        rom[251][38] = 16'h0006;
        rom[251][39] = 16'hFFC0;
        rom[251][40] = 16'h000E;
        rom[251][41] = 16'hFFE6;
        rom[251][42] = 16'h0026;
        rom[251][43] = 16'hFFE0;
        rom[251][44] = 16'h0001;
        rom[251][45] = 16'h0015;
        rom[251][46] = 16'hFFF9;
        rom[251][47] = 16'h002E;
        rom[251][48] = 16'hFFFA;
        rom[251][49] = 16'hFFF9;
        rom[251][50] = 16'h0023;
        rom[251][51] = 16'h0041;
        rom[251][52] = 16'hFFD6;
        rom[251][53] = 16'hFFC4;
        rom[251][54] = 16'h0006;
        rom[251][55] = 16'hFFD7;
        rom[251][56] = 16'h001C;
        rom[251][57] = 16'h000B;
        rom[251][58] = 16'h0008;
        rom[251][59] = 16'h0002;
        rom[251][60] = 16'hFFEF;
        rom[251][61] = 16'h0002;
        rom[251][62] = 16'hFFE0;
        rom[251][63] = 16'h0005;
        rom[251][64] = 16'h0014;
        rom[251][65] = 16'hFFE6;
        rom[251][66] = 16'hFFD7;
        rom[251][67] = 16'h0008;
        rom[251][68] = 16'hFFF1;
        rom[251][69] = 16'hFFDC;
        rom[251][70] = 16'h0005;
        rom[251][71] = 16'h0002;
        rom[251][72] = 16'h002D;
        rom[251][73] = 16'hFFFE;
        rom[251][74] = 16'h0017;
        rom[251][75] = 16'hFFEB;
        rom[251][76] = 16'hFFE2;
        rom[251][77] = 16'h0000;
        rom[251][78] = 16'hFFFE;
        rom[251][79] = 16'h0024;
        rom[251][80] = 16'hFFDC;
        rom[251][81] = 16'h0012;
        rom[251][82] = 16'h000C;
        rom[251][83] = 16'h000D;
        rom[251][84] = 16'hFFEC;
        rom[251][85] = 16'hFFF7;
        rom[251][86] = 16'h0011;
        rom[251][87] = 16'hFFE3;
        rom[251][88] = 16'hFFE8;
        rom[251][89] = 16'h0011;
        rom[251][90] = 16'h0034;
        rom[251][91] = 16'hFFEF;
        rom[251][92] = 16'hFFD9;
        rom[251][93] = 16'h001B;
        rom[251][94] = 16'hFFC9;
        rom[251][95] = 16'hFFE6;
        rom[251][96] = 16'hFFF8;
        rom[251][97] = 16'hFFFE;
        rom[251][98] = 16'h0003;
        rom[251][99] = 16'hFFFC;
        rom[251][100] = 16'hFFFA;
        rom[251][101] = 16'h0000;
        rom[251][102] = 16'h0000;
        rom[251][103] = 16'h0007;
        rom[251][104] = 16'h0015;
        rom[251][105] = 16'hFFEF;
        rom[251][106] = 16'hFFFC;
        rom[251][107] = 16'h0011;
        rom[251][108] = 16'h0011;
        rom[251][109] = 16'h0007;
        rom[251][110] = 16'h0020;
        rom[251][111] = 16'hFFF2;
        rom[251][112] = 16'h0016;
        rom[251][113] = 16'h0017;
        rom[251][114] = 16'hFFFE;
        rom[251][115] = 16'hFFE5;
        rom[251][116] = 16'hFFF4;
        rom[251][117] = 16'hFFC3;
        rom[251][118] = 16'hFFF2;
        rom[251][119] = 16'h002E;
        rom[251][120] = 16'hFFF7;
        rom[251][121] = 16'hFFE0;
        rom[251][122] = 16'h0002;
        rom[251][123] = 16'hFFDE;
        rom[251][124] = 16'hFFF8;
        rom[251][125] = 16'h003D;
        rom[251][126] = 16'hFFF7;
        rom[251][127] = 16'hFFFF;
        rom[252][0] = 16'hFFFE;
        rom[252][1] = 16'hFFAD;
        rom[252][2] = 16'hFFEE;
        rom[252][3] = 16'h001B;
        rom[252][4] = 16'h0012;
        rom[252][5] = 16'hFFF4;
        rom[252][6] = 16'h000C;
        rom[252][7] = 16'hFFC5;
        rom[252][8] = 16'h0023;
        rom[252][9] = 16'hFFE7;
        rom[252][10] = 16'hFFF7;
        rom[252][11] = 16'hFFF0;
        rom[252][12] = 16'h000E;
        rom[252][13] = 16'h000F;
        rom[252][14] = 16'hFFED;
        rom[252][15] = 16'hFFF2;
        rom[252][16] = 16'hFFE1;
        rom[252][17] = 16'hFFCE;
        rom[252][18] = 16'hFFEF;
        rom[252][19] = 16'hFFE3;
        rom[252][20] = 16'hFFFC;
        rom[252][21] = 16'hFFE2;
        rom[252][22] = 16'h0022;
        rom[252][23] = 16'hFFD3;
        rom[252][24] = 16'hFFC8;
        rom[252][25] = 16'h0005;
        rom[252][26] = 16'hFFE6;
        rom[252][27] = 16'h0022;
        rom[252][28] = 16'hFFFC;
        rom[252][29] = 16'hFFF5;
        rom[252][30] = 16'hFFF3;
        rom[252][31] = 16'hFFFB;
        rom[252][32] = 16'h0016;
        rom[252][33] = 16'hFFCA;
        rom[252][34] = 16'h0023;
        rom[252][35] = 16'h0011;
        rom[252][36] = 16'hFFED;
        rom[252][37] = 16'hFFB3;
        rom[252][38] = 16'hFFCC;
        rom[252][39] = 16'h0014;
        rom[252][40] = 16'h001B;
        rom[252][41] = 16'h001A;
        rom[252][42] = 16'hFFF8;
        rom[252][43] = 16'h0003;
        rom[252][44] = 16'h0017;
        rom[252][45] = 16'h0024;
        rom[252][46] = 16'hFFA9;
        rom[252][47] = 16'h0016;
        rom[252][48] = 16'h0003;
        rom[252][49] = 16'h0001;
        rom[252][50] = 16'hFFF4;
        rom[252][51] = 16'hFFF9;
        rom[252][52] = 16'hFFF8;
        rom[252][53] = 16'h0012;
        rom[252][54] = 16'hFFF5;
        rom[252][55] = 16'h0037;
        rom[252][56] = 16'h0005;
        rom[252][57] = 16'h0020;
        rom[252][58] = 16'hFFF4;
        rom[252][59] = 16'hFFD4;
        rom[252][60] = 16'hFFED;
        rom[252][61] = 16'h001B;
        rom[252][62] = 16'hFFF2;
        rom[252][63] = 16'h0021;
        rom[252][64] = 16'h0044;
        rom[252][65] = 16'hFFA6;
        rom[252][66] = 16'hFFEB;
        rom[252][67] = 16'hFFF2;
        rom[252][68] = 16'hFFFD;
        rom[252][69] = 16'hFFF1;
        rom[252][70] = 16'hFFD6;
        rom[252][71] = 16'h0029;
        rom[252][72] = 16'hFFF7;
        rom[252][73] = 16'h0011;
        rom[252][74] = 16'h0010;
        rom[252][75] = 16'hFFF2;
        rom[252][76] = 16'hFF9D;
        rom[252][77] = 16'hFFF1;
        rom[252][78] = 16'hFFFE;
        rom[252][79] = 16'h0013;
        rom[252][80] = 16'hFFC6;
        rom[252][81] = 16'hFFFC;
        rom[252][82] = 16'hFFDD;
        rom[252][83] = 16'h000F;
        rom[252][84] = 16'hFFEB;
        rom[252][85] = 16'hFFF7;
        rom[252][86] = 16'hFFD7;
        rom[252][87] = 16'h0007;
        rom[252][88] = 16'hFFD2;
        rom[252][89] = 16'h0008;
        rom[252][90] = 16'hFFE1;
        rom[252][91] = 16'hFFFE;
        rom[252][92] = 16'hFFC8;
        rom[252][93] = 16'hFFF6;
        rom[252][94] = 16'hFFE5;
        rom[252][95] = 16'hFFFB;
        rom[252][96] = 16'h0011;
        rom[252][97] = 16'hFFFE;
        rom[252][98] = 16'hFFEB;
        rom[252][99] = 16'h001A;
        rom[252][100] = 16'hFFDC;
        rom[252][101] = 16'hFFFE;
        rom[252][102] = 16'h000C;
        rom[252][103] = 16'hFFE4;
        rom[252][104] = 16'h001B;
        rom[252][105] = 16'hFFFA;
        rom[252][106] = 16'hFFDF;
        rom[252][107] = 16'hFFED;
        rom[252][108] = 16'hFFC6;
        rom[252][109] = 16'h000C;
        rom[252][110] = 16'hFFE2;
        rom[252][111] = 16'hFFF8;
        rom[252][112] = 16'hFFE5;
        rom[252][113] = 16'h0031;
        rom[252][114] = 16'hFFF8;
        rom[252][115] = 16'hFFE7;
        rom[252][116] = 16'hFFB0;
        rom[252][117] = 16'hFFE4;
        rom[252][118] = 16'hFFEE;
        rom[252][119] = 16'hFFFA;
        rom[252][120] = 16'hFFDF;
        rom[252][121] = 16'hFFFC;
        rom[252][122] = 16'hFFE8;
        rom[252][123] = 16'hFFAA;
        rom[252][124] = 16'h0008;
        rom[252][125] = 16'h0016;
        rom[252][126] = 16'h0007;
        rom[252][127] = 16'h0016;
        rom[253][0] = 16'hFFE9;
        rom[253][1] = 16'hFFE1;
        rom[253][2] = 16'hFFF5;
        rom[253][3] = 16'h001C;
        rom[253][4] = 16'h001B;
        rom[253][5] = 16'hFFDE;
        rom[253][6] = 16'hFFEE;
        rom[253][7] = 16'hFFD9;
        rom[253][8] = 16'hFFC5;
        rom[253][9] = 16'h0010;
        rom[253][10] = 16'h0000;
        rom[253][11] = 16'hFFDF;
        rom[253][12] = 16'h001D;
        rom[253][13] = 16'hFFD5;
        rom[253][14] = 16'hFFF3;
        rom[253][15] = 16'hFFFE;
        rom[253][16] = 16'h001D;
        rom[253][17] = 16'hFFC2;
        rom[253][18] = 16'h0007;
        rom[253][19] = 16'hFFE3;
        rom[253][20] = 16'hFFF8;
        rom[253][21] = 16'hFFE7;
        rom[253][22] = 16'hFFE9;
        rom[253][23] = 16'hFFBA;
        rom[253][24] = 16'h0003;
        rom[253][25] = 16'hFFDD;
        rom[253][26] = 16'hFFFA;
        rom[253][27] = 16'h0033;
        rom[253][28] = 16'h0010;
        rom[253][29] = 16'hFFB4;
        rom[253][30] = 16'h0007;
        rom[253][31] = 16'hFFED;
        rom[253][32] = 16'hFFFE;
        rom[253][33] = 16'hFFBF;
        rom[253][34] = 16'hFFEC;
        rom[253][35] = 16'h0002;
        rom[253][36] = 16'h001A;
        rom[253][37] = 16'hFFC4;
        rom[253][38] = 16'hFFD6;
        rom[253][39] = 16'hFFD8;
        rom[253][40] = 16'hFFE6;
        rom[253][41] = 16'hFFC7;
        rom[253][42] = 16'h000E;
        rom[253][43] = 16'h0016;
        rom[253][44] = 16'hFFE6;
        rom[253][45] = 16'h000D;
        rom[253][46] = 16'h0008;
        rom[253][47] = 16'h0016;
        rom[253][48] = 16'hFFF7;
        rom[253][49] = 16'h0002;
        rom[253][50] = 16'hFFFE;
        rom[253][51] = 16'hFFF9;
        rom[253][52] = 16'hFFFA;
        rom[253][53] = 16'hFFEB;
        rom[253][54] = 16'h000C;
        rom[253][55] = 16'hFFC0;
        rom[253][56] = 16'hFFE1;
        rom[253][57] = 16'h0007;
        rom[253][58] = 16'h0031;
        rom[253][59] = 16'h0029;
        rom[253][60] = 16'h0006;
        rom[253][61] = 16'h0010;
        rom[253][62] = 16'hFFF9;
        rom[253][63] = 16'hFFA2;
        rom[253][64] = 16'h000F;
        rom[253][65] = 16'h0001;
        rom[253][66] = 16'hFFE1;
        rom[253][67] = 16'hFFDD;
        rom[253][68] = 16'hFFFA;
        rom[253][69] = 16'hFFD7;
        rom[253][70] = 16'hFFEA;
        rom[253][71] = 16'h0007;
        rom[253][72] = 16'h0018;
        rom[253][73] = 16'h0005;
        rom[253][74] = 16'h0005;
        rom[253][75] = 16'hFFC3;
        rom[253][76] = 16'h0022;
        rom[253][77] = 16'h0014;
        rom[253][78] = 16'h000B;
        rom[253][79] = 16'h0038;
        rom[253][80] = 16'hFFD1;
        rom[253][81] = 16'h0008;
        rom[253][82] = 16'hFFCF;
        rom[253][83] = 16'hFFD4;
        rom[253][84] = 16'hFFFA;
        rom[253][85] = 16'h001A;
        rom[253][86] = 16'hFFDC;
        rom[253][87] = 16'h0011;
        rom[253][88] = 16'hFFCF;
        rom[253][89] = 16'h001D;
        rom[253][90] = 16'hFFEB;
        rom[253][91] = 16'h001C;
        rom[253][92] = 16'hFFEB;
        rom[253][93] = 16'hFFE5;
        rom[253][94] = 16'hFFEF;
        rom[253][95] = 16'hFFE2;
        rom[253][96] = 16'h0003;
        rom[253][97] = 16'hFFD0;
        rom[253][98] = 16'h0011;
        rom[253][99] = 16'hFFF1;
        rom[253][100] = 16'h0029;
        rom[253][101] = 16'h0008;
        rom[253][102] = 16'hFFD4;
        rom[253][103] = 16'hFFDD;
        rom[253][104] = 16'h0029;
        rom[253][105] = 16'hFFDD;
        rom[253][106] = 16'h000D;
        rom[253][107] = 16'hFFF0;
        rom[253][108] = 16'hFFFA;
        rom[253][109] = 16'h0015;
        rom[253][110] = 16'hFFEA;
        rom[253][111] = 16'h000A;
        rom[253][112] = 16'hFFFE;
        rom[253][113] = 16'hFF9C;
        rom[253][114] = 16'h0011;
        rom[253][115] = 16'hFFCC;
        rom[253][116] = 16'hFFF3;
        rom[253][117] = 16'hFFE7;
        rom[253][118] = 16'h001D;
        rom[253][119] = 16'h0002;
        rom[253][120] = 16'h0007;
        rom[253][121] = 16'h0002;
        rom[253][122] = 16'h0021;
        rom[253][123] = 16'hFFFE;
        rom[253][124] = 16'h000B;
        rom[253][125] = 16'h0011;
        rom[253][126] = 16'h001A;
        rom[253][127] = 16'h0005;
        rom[254][0] = 16'h0003;
        rom[254][1] = 16'hFFF9;
        rom[254][2] = 16'hFFDF;
        rom[254][3] = 16'hFFE7;
        rom[254][4] = 16'h0040;
        rom[254][5] = 16'hFFF9;
        rom[254][6] = 16'hFFE1;
        rom[254][7] = 16'h001B;
        rom[254][8] = 16'h001E;
        rom[254][9] = 16'h0005;
        rom[254][10] = 16'h000D;
        rom[254][11] = 16'hFFC0;
        rom[254][12] = 16'h0001;
        rom[254][13] = 16'h0013;
        rom[254][14] = 16'hFFCB;
        rom[254][15] = 16'hFFDC;
        rom[254][16] = 16'hFFEF;
        rom[254][17] = 16'h0011;
        rom[254][18] = 16'hFFF1;
        rom[254][19] = 16'h001B;
        rom[254][20] = 16'hFFFC;
        rom[254][21] = 16'h0002;
        rom[254][22] = 16'hFFF1;
        rom[254][23] = 16'hFFE5;
        rom[254][24] = 16'hFFC2;
        rom[254][25] = 16'h0016;
        rom[254][26] = 16'hFFF6;
        rom[254][27] = 16'h0012;
        rom[254][28] = 16'hFFEE;
        rom[254][29] = 16'h0015;
        rom[254][30] = 16'hFFE4;
        rom[254][31] = 16'hFFDC;
        rom[254][32] = 16'h0030;
        rom[254][33] = 16'h0026;
        rom[254][34] = 16'hFFE4;
        rom[254][35] = 16'hFFC8;
        rom[254][36] = 16'h0014;
        rom[254][37] = 16'hFFF8;
        rom[254][38] = 16'h001C;
        rom[254][39] = 16'h000E;
        rom[254][40] = 16'h0024;
        rom[254][41] = 16'hFFF7;
        rom[254][42] = 16'h0007;
        rom[254][43] = 16'h000C;
        rom[254][44] = 16'h000F;
        rom[254][45] = 16'hFFF4;
        rom[254][46] = 16'hFFF9;
        rom[254][47] = 16'h000D;
        rom[254][48] = 16'h0029;
        rom[254][49] = 16'h0023;
        rom[254][50] = 16'hFFEF;
        rom[254][51] = 16'h0023;
        rom[254][52] = 16'h001A;
        rom[254][53] = 16'h0011;
        rom[254][54] = 16'h0006;
        rom[254][55] = 16'hFFFE;
        rom[254][56] = 16'h0016;
        rom[254][57] = 16'h0020;
        rom[254][58] = 16'h001F;
        rom[254][59] = 16'hFFCD;
        rom[254][60] = 16'hFFE5;
        rom[254][61] = 16'h0033;
        rom[254][62] = 16'hFFA5;
        rom[254][63] = 16'hFFF8;
        rom[254][64] = 16'hFFE5;
        rom[254][65] = 16'hFFDB;
        rom[254][66] = 16'hFFF4;
        rom[254][67] = 16'h0044;
        rom[254][68] = 16'h0038;
        rom[254][69] = 16'hFFDB;
        rom[254][70] = 16'hFFF2;
        rom[254][71] = 16'hFFD6;
        rom[254][72] = 16'h000B;
        rom[254][73] = 16'h002C;
        rom[254][74] = 16'h0012;
        rom[254][75] = 16'hFFFE;
        rom[254][76] = 16'hFFDB;
        rom[254][77] = 16'hFFF4;
        rom[254][78] = 16'hFFFE;
        rom[254][79] = 16'h000A;
        rom[254][80] = 16'hFFE2;
        rom[254][81] = 16'hFFE9;
        rom[254][82] = 16'hFFF8;
        rom[254][83] = 16'h001E;
        rom[254][84] = 16'h002C;
        rom[254][85] = 16'hFFF6;
        rom[254][86] = 16'hFFE5;
        rom[254][87] = 16'h000F;
        rom[254][88] = 16'hFFE1;
        rom[254][89] = 16'h000C;
        rom[254][90] = 16'h0019;
        rom[254][91] = 16'hFFCB;
        rom[254][92] = 16'hFFB1;
        rom[254][93] = 16'hFFD7;
        rom[254][94] = 16'h0033;
        rom[254][95] = 16'h0024;
        rom[254][96] = 16'h0009;
        rom[254][97] = 16'h0021;
        rom[254][98] = 16'hFFC3;
        rom[254][99] = 16'hFFDE;
        rom[254][100] = 16'hFFB7;
        rom[254][101] = 16'hFFE2;
        rom[254][102] = 16'hFFF9;
        rom[254][103] = 16'hFFF5;
        rom[254][104] = 16'h0002;
        rom[254][105] = 16'hFFF0;
        rom[254][106] = 16'hFFFB;
        rom[254][107] = 16'hFFE1;
        rom[254][108] = 16'h0009;
        rom[254][109] = 16'hFFFA;
        rom[254][110] = 16'h0022;
        rom[254][111] = 16'hFF9F;
        rom[254][112] = 16'h003F;
        rom[254][113] = 16'h0033;
        rom[254][114] = 16'hFFCE;
        rom[254][115] = 16'hFFF4;
        rom[254][116] = 16'h0010;
        rom[254][117] = 16'hFFF8;
        rom[254][118] = 16'hFFF4;
        rom[254][119] = 16'h0000;
        rom[254][120] = 16'hFFFE;
        rom[254][121] = 16'hFFE1;
        rom[254][122] = 16'hFFD7;
        rom[254][123] = 16'hFFDF;
        rom[254][124] = 16'hFFFD;
        rom[254][125] = 16'h001F;
        rom[254][126] = 16'h0012;
        rom[254][127] = 16'h0047;
        rom[255][0] = 16'hFFDB;
        rom[255][1] = 16'h001D;
        rom[255][2] = 16'h000F;
        rom[255][3] = 16'hFFFD;
        rom[255][4] = 16'hFFD6;
        rom[255][5] = 16'h0010;
        rom[255][6] = 16'hFFFC;
        rom[255][7] = 16'hFFF8;
        rom[255][8] = 16'hFFF1;
        rom[255][9] = 16'h001B;
        rom[255][10] = 16'hFFF9;
        rom[255][11] = 16'hFFE2;
        rom[255][12] = 16'hFFD2;
        rom[255][13] = 16'hFFC9;
        rom[255][14] = 16'hFFC3;
        rom[255][15] = 16'hFFFF;
        rom[255][16] = 16'h0000;
        rom[255][17] = 16'hFFDF;
        rom[255][18] = 16'hFFE2;
        rom[255][19] = 16'h0013;
        rom[255][20] = 16'hFFF4;
        rom[255][21] = 16'h0012;
        rom[255][22] = 16'h001E;
        rom[255][23] = 16'hFFDC;
        rom[255][24] = 16'h0009;
        rom[255][25] = 16'hFFD4;
        rom[255][26] = 16'hFFD1;
        rom[255][27] = 16'hFFF1;
        rom[255][28] = 16'h000D;
        rom[255][29] = 16'hFFFE;
        rom[255][30] = 16'hFFD0;
        rom[255][31] = 16'hFFCD;
        rom[255][32] = 16'h000D;
        rom[255][33] = 16'hFFDC;
        rom[255][34] = 16'hFFD3;
        rom[255][35] = 16'hFFF9;
        rom[255][36] = 16'hFFFA;
        rom[255][37] = 16'hFFDC;
        rom[255][38] = 16'h001A;
        rom[255][39] = 16'hFFF3;
        rom[255][40] = 16'hFFB5;
        rom[255][41] = 16'hFFE5;
        rom[255][42] = 16'hFFDB;
        rom[255][43] = 16'h000D;
        rom[255][44] = 16'hFFD2;
        rom[255][45] = 16'hFFF6;
        rom[255][46] = 16'hFFE9;
        rom[255][47] = 16'hFFD8;
        rom[255][48] = 16'h000A;
        rom[255][49] = 16'h0019;
        rom[255][50] = 16'h000D;
        rom[255][51] = 16'hFFD7;
        rom[255][52] = 16'h000A;
        rom[255][53] = 16'hFFC1;
        rom[255][54] = 16'hFFD9;
        rom[255][55] = 16'hFFE8;
        rom[255][56] = 16'hFFFB;
        rom[255][57] = 16'hFFE5;
        rom[255][58] = 16'h0008;
        rom[255][59] = 16'hFFC2;
        rom[255][60] = 16'h0006;
        rom[255][61] = 16'h001D;
        rom[255][62] = 16'hFFE4;
        rom[255][63] = 16'hFFE8;
        rom[255][64] = 16'h000D;
        rom[255][65] = 16'hFFC6;
        rom[255][66] = 16'hFFEA;
        rom[255][67] = 16'hFFFD;
        rom[255][68] = 16'hFFDF;
        rom[255][69] = 16'hFFFE;
        rom[255][70] = 16'h0014;
        rom[255][71] = 16'hFFFA;
        rom[255][72] = 16'hFFBD;
        rom[255][73] = 16'hFFF8;
        rom[255][74] = 16'hFFD1;
        rom[255][75] = 16'hFFFC;
        rom[255][76] = 16'h0007;
        rom[255][77] = 16'hFFD2;
        rom[255][78] = 16'hFFEF;
        rom[255][79] = 16'hFFE6;
        rom[255][80] = 16'hFFF8;
        rom[255][81] = 16'h001A;
        rom[255][82] = 16'h0003;
        rom[255][83] = 16'hFFF4;
        rom[255][84] = 16'h0019;
        rom[255][85] = 16'hFFF9;
        rom[255][86] = 16'h000A;
        rom[255][87] = 16'h0011;
        rom[255][88] = 16'hFFD8;
        rom[255][89] = 16'hFFEF;
        rom[255][90] = 16'hFFF3;
        rom[255][91] = 16'h000C;
        rom[255][92] = 16'hFFE5;
        rom[255][93] = 16'hFFF5;
        rom[255][94] = 16'hFFC9;
        rom[255][95] = 16'hFFF3;
        rom[255][96] = 16'h000A;
        rom[255][97] = 16'hFFFF;
        rom[255][98] = 16'hFFF4;
        rom[255][99] = 16'h000F;
        rom[255][100] = 16'hFFF4;
        rom[255][101] = 16'hFFD9;
        rom[255][102] = 16'hFFFE;
        rom[255][103] = 16'h0007;
        rom[255][104] = 16'hFFCB;
        rom[255][105] = 16'hFFF2;
        rom[255][106] = 16'h0002;
        rom[255][107] = 16'hFFEF;
        rom[255][108] = 16'h000C;
        rom[255][109] = 16'h001E;
        rom[255][110] = 16'hFFE7;
        rom[255][111] = 16'h0015;
        rom[255][112] = 16'hFFF2;
        rom[255][113] = 16'h0011;
        rom[255][114] = 16'hFFEF;
        rom[255][115] = 16'hFFB2;
        rom[255][116] = 16'hFFF5;
        rom[255][117] = 16'hFFED;
        rom[255][118] = 16'hFFD0;
        rom[255][119] = 16'h0004;
        rom[255][120] = 16'hFFBE;
        rom[255][121] = 16'hFFF1;
        rom[255][122] = 16'hFFD9;
        rom[255][123] = 16'h0007;
        rom[255][124] = 16'hFFFF;
        rom[255][125] = 16'hFFCD;
        rom[255][126] = 16'hFFE4;
        rom[255][127] = 16'hFFEF;
    end

    always @(*) begin
        data_out = rom[addr][index];
    end
endmodule
