// Q8.8 Fixed-Point ROM: rom_layer4_weights
module rom_layer4_weights (
    input [6:0] addr,
    input [3:0] index,
    output reg signed [15:0] data_out
);

    reg signed [15:0] rom [0:127][0:9];

    initial begin
        rom[0][0] = 16'h0037;
        rom[0][1] = 16'h0027;
        rom[0][2] = 16'hFFC3;
        rom[0][3] = 16'h0012;
        rom[0][4] = 16'h0037;
        rom[0][5] = 16'h002C;
        rom[0][6] = 16'h0037;
        rom[0][7] = 16'hFFC6;
        rom[0][8] = 16'hFFE3;
        rom[0][9] = 16'h0031;
        rom[1][0] = 16'h0001;
        rom[1][1] = 16'h0022;
        rom[1][2] = 16'h000F;
        rom[1][3] = 16'hFFFA;
        rom[1][4] = 16'hFFF2;
        rom[1][5] = 16'hFFFA;
        rom[1][6] = 16'hFFE1;
        rom[1][7] = 16'h002C;
        rom[1][8] = 16'h002F;
        rom[1][9] = 16'hFFDD;
        rom[2][0] = 16'hFFE7;
        rom[2][1] = 16'hFFD3;
        rom[2][2] = 16'hFFC9;
        rom[2][3] = 16'h0015;
        rom[2][4] = 16'hFFD6;
        rom[2][5] = 16'h0017;
        rom[2][6] = 16'h0017;
        rom[2][7] = 16'hFFDC;
        rom[2][8] = 16'hFFED;
        rom[2][9] = 16'h0011;
        rom[3][0] = 16'hFFBD;
        rom[3][1] = 16'h000C;
        rom[3][2] = 16'hFFE1;
        rom[3][3] = 16'h0014;
        rom[3][4] = 16'hFFE6;
        rom[3][5] = 16'hFFE2;
        rom[3][6] = 16'hFFE8;
        rom[3][7] = 16'h0040;
        rom[3][8] = 16'hFFC3;
        rom[3][9] = 16'h002B;
        rom[4][0] = 16'hFFF1;
        rom[4][1] = 16'hFFD4;
        rom[4][2] = 16'hFFE5;
        rom[4][3] = 16'hFFC5;
        rom[4][4] = 16'h000F;
        rom[4][5] = 16'hFFBF;
        rom[4][6] = 16'hFFE9;
        rom[4][7] = 16'hFFF1;
        rom[4][8] = 16'h0015;
        rom[4][9] = 16'hFFCE;
        rom[5][0] = 16'h0006;
        rom[5][1] = 16'hFFEF;
        rom[5][2] = 16'hFFE9;
        rom[5][3] = 16'h000E;
        rom[5][4] = 16'h002D;
        rom[5][5] = 16'h0006;
        rom[5][6] = 16'hFFF1;
        rom[5][7] = 16'h0035;
        rom[5][8] = 16'h003A;
        rom[5][9] = 16'hFFD8;
        rom[6][0] = 16'h0029;
        rom[6][1] = 16'h0030;
        rom[6][2] = 16'h003E;
        rom[6][3] = 16'hFFDD;
        rom[6][4] = 16'hFFDD;
        rom[6][5] = 16'hFFEE;
        rom[6][6] = 16'hFFD7;
        rom[6][7] = 16'h003B;
        rom[6][8] = 16'h000D;
        rom[6][9] = 16'h0030;
        rom[7][0] = 16'h0020;
        rom[7][1] = 16'h001D;
        rom[7][2] = 16'h002F;
        rom[7][3] = 16'h0000;
        rom[7][4] = 16'hFFB2;
        rom[7][5] = 16'hFFE9;
        rom[7][6] = 16'hFFCB;
        rom[7][7] = 16'h001D;
        rom[7][8] = 16'h000E;
        rom[7][9] = 16'hFFC0;
        rom[8][0] = 16'h0049;
        rom[8][1] = 16'h0017;
        rom[8][2] = 16'hFFF0;
        rom[8][3] = 16'hFFEE;
        rom[8][4] = 16'h0019;
        rom[8][5] = 16'hFFEF;
        rom[8][6] = 16'h0027;
        rom[8][7] = 16'hFFE5;
        rom[8][8] = 16'h0034;
        rom[8][9] = 16'hFFC4;
        rom[9][0] = 16'hFFA3;
        rom[9][1] = 16'h0035;
        rom[9][2] = 16'hFFEE;
        rom[9][3] = 16'h003A;
        rom[9][4] = 16'hFFEB;
        rom[9][5] = 16'h0033;
        rom[9][6] = 16'h001D;
        rom[9][7] = 16'h001B;
        rom[9][8] = 16'hFFCF;
        rom[9][9] = 16'hFFCC;
        rom[10][0] = 16'h000B;
        rom[10][1] = 16'h0029;
        rom[10][2] = 16'h0048;
        rom[10][3] = 16'hFFC6;
        rom[10][4] = 16'hFFBD;
        rom[10][5] = 16'hFFE7;
        rom[10][6] = 16'h0017;
        rom[10][7] = 16'h0011;
        rom[10][8] = 16'hFFD5;
        rom[10][9] = 16'hFFFA;
        rom[11][0] = 16'hFFB4;
        rom[11][1] = 16'hFFE2;
        rom[11][2] = 16'hFFFB;
        rom[11][3] = 16'hFFE8;
        rom[11][4] = 16'h002E;
        rom[11][5] = 16'hFFEA;
        rom[11][6] = 16'h0039;
        rom[11][7] = 16'hFFB2;
        rom[11][8] = 16'hFFDD;
        rom[11][9] = 16'h0015;
        rom[12][0] = 16'hFFD3;
        rom[12][1] = 16'hFFEE;
        rom[12][2] = 16'hFFCA;
        rom[12][3] = 16'h0019;
        rom[12][4] = 16'hFFBF;
        rom[12][5] = 16'hFFE0;
        rom[12][6] = 16'h0032;
        rom[12][7] = 16'hFFDB;
        rom[12][8] = 16'h0000;
        rom[12][9] = 16'hFFC9;
        rom[13][0] = 16'h003E;
        rom[13][1] = 16'hFFE8;
        rom[13][2] = 16'h002B;
        rom[13][3] = 16'h001B;
        rom[13][4] = 16'h001C;
        rom[13][5] = 16'hFFDD;
        rom[13][6] = 16'h000B;
        rom[13][7] = 16'hFFF1;
        rom[13][8] = 16'hFFE9;
        rom[13][9] = 16'h0001;
        rom[14][0] = 16'h0000;
        rom[14][1] = 16'h0018;
        rom[14][2] = 16'h0003;
        rom[14][3] = 16'hFFF3;
        rom[14][4] = 16'hFFBC;
        rom[14][5] = 16'hFFFB;
        rom[14][6] = 16'hFFD9;
        rom[14][7] = 16'h0016;
        rom[14][8] = 16'h0025;
        rom[14][9] = 16'hFF95;
        rom[15][0] = 16'hFFF1;
        rom[15][1] = 16'hFFFD;
        rom[15][2] = 16'hFFD9;
        rom[15][3] = 16'h0008;
        rom[15][4] = 16'hFFF1;
        rom[15][5] = 16'h0009;
        rom[15][6] = 16'hFFCB;
        rom[15][7] = 16'hFFDE;
        rom[15][8] = 16'hFFFA;
        rom[15][9] = 16'hFFF9;
        rom[16][0] = 16'h0008;
        rom[16][1] = 16'h0024;
        rom[16][2] = 16'hFFFD;
        rom[16][3] = 16'h000A;
        rom[16][4] = 16'h001A;
        rom[16][5] = 16'hFFE1;
        rom[16][6] = 16'h0004;
        rom[16][7] = 16'h001D;
        rom[16][8] = 16'hFFC7;
        rom[16][9] = 16'h001B;
        rom[17][0] = 16'h002D;
        rom[17][1] = 16'h000F;
        rom[17][2] = 16'h003D;
        rom[17][3] = 16'h000D;
        rom[17][4] = 16'hFFB4;
        rom[17][5] = 16'hFFD9;
        rom[17][6] = 16'hFFC8;
        rom[17][7] = 16'h0029;
        rom[17][8] = 16'h002F;
        rom[17][9] = 16'hFFC9;
        rom[18][0] = 16'hFFD7;
        rom[18][1] = 16'h0027;
        rom[18][2] = 16'hFFC4;
        rom[18][3] = 16'h0008;
        rom[18][4] = 16'h000D;
        rom[18][5] = 16'hFFFC;
        rom[18][6] = 16'h003C;
        rom[18][7] = 16'hFFF3;
        rom[18][8] = 16'hFFFD;
        rom[18][9] = 16'hFFFA;
        rom[19][0] = 16'h0012;
        rom[19][1] = 16'h002A;
        rom[19][2] = 16'hFFE9;
        rom[19][3] = 16'h0022;
        rom[19][4] = 16'hFFC4;
        rom[19][5] = 16'hFFF5;
        rom[19][6] = 16'hFFBE;
        rom[19][7] = 16'h0018;
        rom[19][8] = 16'h0032;
        rom[19][9] = 16'hFFCE;
        rom[20][0] = 16'hFFB9;
        rom[20][1] = 16'hFFD7;
        rom[20][2] = 16'h0021;
        rom[20][3] = 16'hFFC8;
        rom[20][4] = 16'h0022;
        rom[20][5] = 16'hFFD4;
        rom[20][6] = 16'h002E;
        rom[20][7] = 16'hFFE0;
        rom[20][8] = 16'h0027;
        rom[20][9] = 16'hFFDE;
        rom[21][0] = 16'h0028;
        rom[21][1] = 16'h0011;
        rom[21][2] = 16'hFFFF;
        rom[21][3] = 16'hFFF9;
        rom[21][4] = 16'hFFD4;
        rom[21][5] = 16'h001A;
        rom[21][6] = 16'hFFE3;
        rom[21][7] = 16'hFFE0;
        rom[21][8] = 16'h000F;
        rom[21][9] = 16'hFFF3;
        rom[22][0] = 16'hFFD4;
        rom[22][1] = 16'h0012;
        rom[22][2] = 16'hFFC7;
        rom[22][3] = 16'h0028;
        rom[22][4] = 16'hFFD5;
        rom[22][5] = 16'hFFE2;
        rom[22][6] = 16'hFFDD;
        rom[22][7] = 16'hFFDF;
        rom[22][8] = 16'hFFED;
        rom[22][9] = 16'h0037;
        rom[23][0] = 16'h0016;
        rom[23][1] = 16'h0021;
        rom[23][2] = 16'hFFB6;
        rom[23][3] = 16'hFFB7;
        rom[23][4] = 16'h0032;
        rom[23][5] = 16'hFFBA;
        rom[23][6] = 16'hFFF3;
        rom[23][7] = 16'h0036;
        rom[23][8] = 16'hFFCE;
        rom[23][9] = 16'hFFF8;
        rom[24][0] = 16'hFFF8;
        rom[24][1] = 16'h0006;
        rom[24][2] = 16'hFFC9;
        rom[24][3] = 16'h0005;
        rom[24][4] = 16'hFFEF;
        rom[24][5] = 16'h0016;
        rom[24][6] = 16'hFFC4;
        rom[24][7] = 16'hFFDB;
        rom[24][8] = 16'hFFC4;
        rom[24][9] = 16'hFFC6;
        rom[25][0] = 16'h000A;
        rom[25][1] = 16'hFFD1;
        rom[25][2] = 16'h0027;
        rom[25][3] = 16'hFFC3;
        rom[25][4] = 16'h0015;
        rom[25][5] = 16'hFFB1;
        rom[25][6] = 16'h001B;
        rom[25][7] = 16'h0003;
        rom[25][8] = 16'h001E;
        rom[25][9] = 16'hFF9B;
        rom[26][0] = 16'h0000;
        rom[26][1] = 16'h000A;
        rom[26][2] = 16'h0008;
        rom[26][3] = 16'hFFBF;
        rom[26][4] = 16'hFFF9;
        rom[26][5] = 16'hFFE6;
        rom[26][6] = 16'h001C;
        rom[26][7] = 16'h0003;
        rom[26][8] = 16'h0031;
        rom[26][9] = 16'hFFF9;
        rom[27][0] = 16'hFFAC;
        rom[27][1] = 16'hFFBD;
        rom[27][2] = 16'h0032;
        rom[27][3] = 16'hFFE9;
        rom[27][4] = 16'hFFE2;
        rom[27][5] = 16'hFF9D;
        rom[27][6] = 16'hFFE1;
        rom[27][7] = 16'h0029;
        rom[27][8] = 16'hFFE7;
        rom[27][9] = 16'hFFCF;
        rom[28][0] = 16'hFFD3;
        rom[28][1] = 16'hFFF7;
        rom[28][2] = 16'h0001;
        rom[28][3] = 16'h0020;
        rom[28][4] = 16'hFFC8;
        rom[28][5] = 16'h0017;
        rom[28][6] = 16'hFF9A;
        rom[28][7] = 16'h0020;
        rom[28][8] = 16'h0009;
        rom[28][9] = 16'hFFF2;
        rom[29][0] = 16'h0004;
        rom[29][1] = 16'h0008;
        rom[29][2] = 16'h0031;
        rom[29][3] = 16'h0037;
        rom[29][4] = 16'hFFC9;
        rom[29][5] = 16'h0020;
        rom[29][6] = 16'hFFF0;
        rom[29][7] = 16'hFFEB;
        rom[29][8] = 16'h0024;
        rom[29][9] = 16'hFFCF;
        rom[30][0] = 16'h0022;
        rom[30][1] = 16'hFFEA;
        rom[30][2] = 16'hFFF0;
        rom[30][3] = 16'hFFC3;
        rom[30][4] = 16'h0016;
        rom[30][5] = 16'hFFE1;
        rom[30][6] = 16'h0024;
        rom[30][7] = 16'h0001;
        rom[30][8] = 16'h0008;
        rom[30][9] = 16'hFFCA;
        rom[31][0] = 16'h0042;
        rom[31][1] = 16'hFFF8;
        rom[31][2] = 16'h0035;
        rom[31][3] = 16'hFFF9;
        rom[31][4] = 16'hFFE2;
        rom[31][5] = 16'hFFFE;
        rom[31][6] = 16'h0045;
        rom[31][7] = 16'hFFB2;
        rom[31][8] = 16'hFFCC;
        rom[31][9] = 16'hFFD4;
        rom[32][0] = 16'hFFF1;
        rom[32][1] = 16'hFFE3;
        rom[32][2] = 16'hFFD4;
        rom[32][3] = 16'h001F;
        rom[32][4] = 16'hFFD0;
        rom[32][5] = 16'hFFD9;
        rom[32][6] = 16'h0045;
        rom[32][7] = 16'hFFF5;
        rom[32][8] = 16'h001D;
        rom[32][9] = 16'h0019;
        rom[33][0] = 16'h0032;
        rom[33][1] = 16'h0031;
        rom[33][2] = 16'h0024;
        rom[33][3] = 16'hFFF7;
        rom[33][4] = 16'hFFE3;
        rom[33][5] = 16'hFFF8;
        rom[33][6] = 16'hFFB0;
        rom[33][7] = 16'hFFCC;
        rom[33][8] = 16'hFFE0;
        rom[33][9] = 16'hFFF0;
        rom[34][0] = 16'h0043;
        rom[34][1] = 16'hFFEE;
        rom[34][2] = 16'h0040;
        rom[34][3] = 16'hFFFD;
        rom[34][4] = 16'h0025;
        rom[34][5] = 16'hFFE8;
        rom[34][6] = 16'hFFF9;
        rom[34][7] = 16'hFFEB;
        rom[34][8] = 16'hFFC9;
        rom[34][9] = 16'h003A;
        rom[35][0] = 16'h0012;
        rom[35][1] = 16'hFFDA;
        rom[35][2] = 16'h002B;
        rom[35][3] = 16'h002B;
        rom[35][4] = 16'hFFD9;
        rom[35][5] = 16'h0022;
        rom[35][6] = 16'hFFEB;
        rom[35][7] = 16'hFFF3;
        rom[35][8] = 16'hFFD8;
        rom[35][9] = 16'hFFFA;
        rom[36][0] = 16'h0016;
        rom[36][1] = 16'h001F;
        rom[36][2] = 16'h0022;
        rom[36][3] = 16'h0008;
        rom[36][4] = 16'hFFCB;
        rom[36][5] = 16'hFFCB;
        rom[36][6] = 16'hFFDE;
        rom[36][7] = 16'h001E;
        rom[36][8] = 16'hFFFF;
        rom[36][9] = 16'hFFD8;
        rom[37][0] = 16'hFFDA;
        rom[37][1] = 16'h0008;
        rom[37][2] = 16'hFFDA;
        rom[37][3] = 16'hFFDB;
        rom[37][4] = 16'h0026;
        rom[37][5] = 16'h002B;
        rom[37][6] = 16'hFFE3;
        rom[37][7] = 16'hFFF5;
        rom[37][8] = 16'h002D;
        rom[37][9] = 16'hFFE7;
        rom[38][0] = 16'h0005;
        rom[38][1] = 16'h0037;
        rom[38][2] = 16'hFFCD;
        rom[38][3] = 16'h0036;
        rom[38][4] = 16'hFFEA;
        rom[38][5] = 16'h0033;
        rom[38][6] = 16'hFFAF;
        rom[38][7] = 16'h0024;
        rom[38][8] = 16'hFFC4;
        rom[38][9] = 16'hFFCC;
        rom[39][0] = 16'h004A;
        rom[39][1] = 16'h0032;
        rom[39][2] = 16'h002B;
        rom[39][3] = 16'h0031;
        rom[39][4] = 16'h001B;
        rom[39][5] = 16'h0033;
        rom[39][6] = 16'h0011;
        rom[39][7] = 16'hFFF4;
        rom[39][8] = 16'hFFE5;
        rom[39][9] = 16'h0003;
        rom[40][0] = 16'hFFD9;
        rom[40][1] = 16'hFFB8;
        rom[40][2] = 16'h002F;
        rom[40][3] = 16'h0051;
        rom[40][4] = 16'h0004;
        rom[40][5] = 16'hFFF3;
        rom[40][6] = 16'h0017;
        rom[40][7] = 16'hFFE9;
        rom[40][8] = 16'hFFE7;
        rom[40][9] = 16'hFFE8;
        rom[41][0] = 16'h0020;
        rom[41][1] = 16'h0031;
        rom[41][2] = 16'hFFDC;
        rom[41][3] = 16'h0003;
        rom[41][4] = 16'hFFE4;
        rom[41][5] = 16'h002F;
        rom[41][6] = 16'hFFFD;
        rom[41][7] = 16'hFFD0;
        rom[41][8] = 16'h0001;
        rom[41][9] = 16'hFFCC;
        rom[42][0] = 16'h0002;
        rom[42][1] = 16'hFFFE;
        rom[42][2] = 16'h001D;
        rom[42][3] = 16'hFFE6;
        rom[42][4] = 16'hFFD9;
        rom[42][5] = 16'hFFC8;
        rom[42][6] = 16'h002C;
        rom[42][7] = 16'hFFCB;
        rom[42][8] = 16'hFFE7;
        rom[42][9] = 16'h0051;
        rom[43][0] = 16'hFFCC;
        rom[43][1] = 16'h0024;
        rom[43][2] = 16'hFFB5;
        rom[43][3] = 16'hFFE3;
        rom[43][4] = 16'hFFC2;
        rom[43][5] = 16'h0008;
        rom[43][6] = 16'h0021;
        rom[43][7] = 16'hFFFA;
        rom[43][8] = 16'hFFA4;
        rom[43][9] = 16'h001B;
        rom[44][0] = 16'h0018;
        rom[44][1] = 16'h0007;
        rom[44][2] = 16'h000C;
        rom[44][3] = 16'h000D;
        rom[44][4] = 16'h000B;
        rom[44][5] = 16'h0002;
        rom[44][6] = 16'h0011;
        rom[44][7] = 16'hFFB2;
        rom[44][8] = 16'hFFBF;
        rom[44][9] = 16'hFFFF;
        rom[45][0] = 16'hFFEE;
        rom[45][1] = 16'hFFF5;
        rom[45][2] = 16'h0006;
        rom[45][3] = 16'h0025;
        rom[45][4] = 16'hFFE9;
        rom[45][5] = 16'h002B;
        rom[45][6] = 16'hFFE0;
        rom[45][7] = 16'hFFDF;
        rom[45][8] = 16'hFFDD;
        rom[45][9] = 16'h002B;
        rom[46][0] = 16'hFFCB;
        rom[46][1] = 16'h001F;
        rom[46][2] = 16'hFFD4;
        rom[46][3] = 16'hFFF3;
        rom[46][4] = 16'h0003;
        rom[46][5] = 16'hFFF8;
        rom[46][6] = 16'h000D;
        rom[46][7] = 16'h0022;
        rom[46][8] = 16'hFFCF;
        rom[46][9] = 16'hFFD2;
        rom[47][0] = 16'hFFDE;
        rom[47][1] = 16'hFFF2;
        rom[47][2] = 16'h001D;
        rom[47][3] = 16'h0012;
        rom[47][4] = 16'hFFCD;
        rom[47][5] = 16'h0012;
        rom[47][6] = 16'h003C;
        rom[47][7] = 16'h001E;
        rom[47][8] = 16'h003E;
        rom[47][9] = 16'hFFF6;
        rom[48][0] = 16'hFFCC;
        rom[48][1] = 16'hFFEF;
        rom[48][2] = 16'h0011;
        rom[48][3] = 16'h0022;
        rom[48][4] = 16'h0002;
        rom[48][5] = 16'hFFE9;
        rom[48][6] = 16'hFFC7;
        rom[48][7] = 16'h0035;
        rom[48][8] = 16'hFFE3;
        rom[48][9] = 16'hFFD3;
        rom[49][0] = 16'hFFC7;
        rom[49][1] = 16'h0000;
        rom[49][2] = 16'h003A;
        rom[49][3] = 16'h001D;
        rom[49][4] = 16'h0021;
        rom[49][5] = 16'hFFF3;
        rom[49][6] = 16'hFFF3;
        rom[49][7] = 16'h0031;
        rom[49][8] = 16'h002D;
        rom[49][9] = 16'hFFCE;
        rom[50][0] = 16'hFFC6;
        rom[50][1] = 16'hFFF5;
        rom[50][2] = 16'hFFA2;
        rom[50][3] = 16'h0013;
        rom[50][4] = 16'hFFE6;
        rom[50][5] = 16'h0014;
        rom[50][6] = 16'hFFD3;
        rom[50][7] = 16'h0017;
        rom[50][8] = 16'hFFDE;
        rom[50][9] = 16'h0012;
        rom[51][0] = 16'h002B;
        rom[51][1] = 16'h0015;
        rom[51][2] = 16'hFFEA;
        rom[51][3] = 16'hFFDE;
        rom[51][4] = 16'h0044;
        rom[51][5] = 16'hFFE8;
        rom[51][6] = 16'h0041;
        rom[51][7] = 16'hFFEE;
        rom[51][8] = 16'hFFE2;
        rom[51][9] = 16'h0030;
        rom[52][0] = 16'hFFBE;
        rom[52][1] = 16'hFFE7;
        rom[52][2] = 16'hFFE6;
        rom[52][3] = 16'hFFDC;
        rom[52][4] = 16'hFFD7;
        rom[52][5] = 16'hFFE4;
        rom[52][6] = 16'hFFEE;
        rom[52][7] = 16'hFFC4;
        rom[52][8] = 16'h0008;
        rom[52][9] = 16'h0020;
        rom[53][0] = 16'hFFC3;
        rom[53][1] = 16'hFFBD;
        rom[53][2] = 16'h001A;
        rom[53][3] = 16'h0026;
        rom[53][4] = 16'h0020;
        rom[53][5] = 16'hFFE8;
        rom[53][6] = 16'hFFED;
        rom[53][7] = 16'hFFD9;
        rom[53][8] = 16'hFFF6;
        rom[53][9] = 16'h0039;
        rom[54][0] = 16'h0016;
        rom[54][1] = 16'h0028;
        rom[54][2] = 16'hFFEA;
        rom[54][3] = 16'hFFF0;
        rom[54][4] = 16'h0015;
        rom[54][5] = 16'h0036;
        rom[54][6] = 16'hFFBF;
        rom[54][7] = 16'hFFEE;
        rom[54][8] = 16'hFFEB;
        rom[54][9] = 16'h0017;
        rom[55][0] = 16'h0032;
        rom[55][1] = 16'hFFBE;
        rom[55][2] = 16'h002E;
        rom[55][3] = 16'hFFEF;
        rom[55][4] = 16'hFFE8;
        rom[55][5] = 16'hFFF4;
        rom[55][6] = 16'hFFED;
        rom[55][7] = 16'hFFDD;
        rom[55][8] = 16'h0021;
        rom[55][9] = 16'hFFF7;
        rom[56][0] = 16'h000D;
        rom[56][1] = 16'hFFEF;
        rom[56][2] = 16'h0021;
        rom[56][3] = 16'h0018;
        rom[56][4] = 16'h0013;
        rom[56][5] = 16'h0014;
        rom[56][6] = 16'h001E;
        rom[56][7] = 16'hFFC7;
        rom[56][8] = 16'h001D;
        rom[56][9] = 16'hFFDA;
        rom[57][0] = 16'h003C;
        rom[57][1] = 16'hFFE1;
        rom[57][2] = 16'hFFAA;
        rom[57][3] = 16'hFFD7;
        rom[57][4] = 16'h002D;
        rom[57][5] = 16'hFFC5;
        rom[57][6] = 16'h001D;
        rom[57][7] = 16'h0016;
        rom[57][8] = 16'hFFD6;
        rom[57][9] = 16'h000F;
        rom[58][0] = 16'hFFD3;
        rom[58][1] = 16'hFFFE;
        rom[58][2] = 16'h000D;
        rom[58][3] = 16'hFFC5;
        rom[58][4] = 16'hFFEE;
        rom[58][5] = 16'hFFF3;
        rom[58][6] = 16'h0012;
        rom[58][7] = 16'hFFF3;
        rom[58][8] = 16'hFFCE;
        rom[58][9] = 16'hFFCD;
        rom[59][0] = 16'hFFBA;
        rom[59][1] = 16'hFFF4;
        rom[59][2] = 16'h0017;
        rom[59][3] = 16'hFFDB;
        rom[59][4] = 16'h001A;
        rom[59][5] = 16'hFFE3;
        rom[59][6] = 16'h0027;
        rom[59][7] = 16'h0020;
        rom[59][8] = 16'h001C;
        rom[59][9] = 16'hFFDB;
        rom[60][0] = 16'h0032;
        rom[60][1] = 16'h0015;
        rom[60][2] = 16'hFFB5;
        rom[60][3] = 16'h0013;
        rom[60][4] = 16'h0024;
        rom[60][5] = 16'hFFF1;
        rom[60][6] = 16'hFFFA;
        rom[60][7] = 16'hFFDC;
        rom[60][8] = 16'hFFF5;
        rom[60][9] = 16'hFFEA;
        rom[61][0] = 16'h0007;
        rom[61][1] = 16'hFFEB;
        rom[61][2] = 16'h002C;
        rom[61][3] = 16'h002C;
        rom[61][4] = 16'hFFC9;
        rom[61][5] = 16'hFFF0;
        rom[61][6] = 16'h0020;
        rom[61][7] = 16'hFFE9;
        rom[61][8] = 16'h0016;
        rom[61][9] = 16'hFFD4;
        rom[62][0] = 16'hFFDC;
        rom[62][1] = 16'h0002;
        rom[62][2] = 16'h0014;
        rom[62][3] = 16'hFFF2;
        rom[62][4] = 16'hFFB7;
        rom[62][5] = 16'h0003;
        rom[62][6] = 16'hFFAC;
        rom[62][7] = 16'h000E;
        rom[62][8] = 16'h000D;
        rom[62][9] = 16'hFFB6;
        rom[63][0] = 16'h0012;
        rom[63][1] = 16'hFFE1;
        rom[63][2] = 16'h002B;
        rom[63][3] = 16'hFFC0;
        rom[63][4] = 16'h0000;
        rom[63][5] = 16'hFFEC;
        rom[63][6] = 16'h0021;
        rom[63][7] = 16'h0033;
        rom[63][8] = 16'h0005;
        rom[63][9] = 16'hFFFD;
        rom[64][0] = 16'hFFFC;
        rom[64][1] = 16'hFFED;
        rom[64][2] = 16'hFFEE;
        rom[64][3] = 16'h0044;
        rom[64][4] = 16'h0012;
        rom[64][5] = 16'h0034;
        rom[64][6] = 16'h0033;
        rom[64][7] = 16'hFFDF;
        rom[64][8] = 16'h0002;
        rom[64][9] = 16'h0036;
        rom[65][0] = 16'h0039;
        rom[65][1] = 16'h0026;
        rom[65][2] = 16'h0031;
        rom[65][3] = 16'hFFE9;
        rom[65][4] = 16'h0013;
        rom[65][5] = 16'hFFCA;
        rom[65][6] = 16'hFFDF;
        rom[65][7] = 16'h0001;
        rom[65][8] = 16'hFFF8;
        rom[65][9] = 16'h0008;
        rom[66][0] = 16'hFFD6;
        rom[66][1] = 16'hFFE5;
        rom[66][2] = 16'hFFCB;
        rom[66][3] = 16'hFFF3;
        rom[66][4] = 16'h0016;
        rom[66][5] = 16'h0016;
        rom[66][6] = 16'hFFE1;
        rom[66][7] = 16'h0004;
        rom[66][8] = 16'h0033;
        rom[66][9] = 16'h0002;
        rom[67][0] = 16'hFFF1;
        rom[67][1] = 16'hFFF8;
        rom[67][2] = 16'hFFC8;
        rom[67][3] = 16'hFFEE;
        rom[67][4] = 16'h002A;
        rom[67][5] = 16'hFFD9;
        rom[67][6] = 16'h0025;
        rom[67][7] = 16'h0004;
        rom[67][8] = 16'h0031;
        rom[67][9] = 16'h0013;
        rom[68][0] = 16'hFFB4;
        rom[68][1] = 16'hFFF5;
        rom[68][2] = 16'h001F;
        rom[68][3] = 16'hFFE3;
        rom[68][4] = 16'h002A;
        rom[68][5] = 16'h0003;
        rom[68][6] = 16'hFFE8;
        rom[68][7] = 16'hFFC2;
        rom[68][8] = 16'hFFD8;
        rom[68][9] = 16'hFFF3;
        rom[69][0] = 16'h0021;
        rom[69][1] = 16'h0011;
        rom[69][2] = 16'h0011;
        rom[69][3] = 16'h0016;
        rom[69][4] = 16'hFFEA;
        rom[69][5] = 16'hFFD6;
        rom[69][6] = 16'hFFDD;
        rom[69][7] = 16'hFFDE;
        rom[69][8] = 16'h0044;
        rom[69][9] = 16'h0017;
        rom[70][0] = 16'h0011;
        rom[70][1] = 16'h0013;
        rom[70][2] = 16'hFFDD;
        rom[70][3] = 16'h0022;
        rom[70][4] = 16'hFFAB;
        rom[70][5] = 16'h001D;
        rom[70][6] = 16'hFFC2;
        rom[70][7] = 16'h0005;
        rom[70][8] = 16'h0012;
        rom[70][9] = 16'hFFDA;
        rom[71][0] = 16'hFFD4;
        rom[71][1] = 16'hFFE4;
        rom[71][2] = 16'hFFC0;
        rom[71][3] = 16'hFFCE;
        rom[71][4] = 16'hFFF3;
        rom[71][5] = 16'h0005;
        rom[71][6] = 16'h000A;
        rom[71][7] = 16'hFFF3;
        rom[71][8] = 16'hFFB5;
        rom[71][9] = 16'h0032;
        rom[72][0] = 16'h0041;
        rom[72][1] = 16'hFFEB;
        rom[72][2] = 16'hFFEA;
        rom[72][3] = 16'hFFF3;
        rom[72][4] = 16'h0017;
        rom[72][5] = 16'h000B;
        rom[72][6] = 16'h002E;
        rom[72][7] = 16'hFFCE;
        rom[72][8] = 16'h000D;
        rom[72][9] = 16'hFFD4;
        rom[73][0] = 16'hFFEC;
        rom[73][1] = 16'h0003;
        rom[73][2] = 16'h000E;
        rom[73][3] = 16'h0019;
        rom[73][4] = 16'h001E;
        rom[73][5] = 16'h0016;
        rom[73][6] = 16'h0017;
        rom[73][7] = 16'hFFEF;
        rom[73][8] = 16'h0030;
        rom[73][9] = 16'hFFE9;
        rom[74][0] = 16'h0024;
        rom[74][1] = 16'hFFCC;
        rom[74][2] = 16'h0043;
        rom[74][3] = 16'hFFE6;
        rom[74][4] = 16'hFFFE;
        rom[74][5] = 16'hFFF7;
        rom[74][6] = 16'h002B;
        rom[74][7] = 16'hFFF0;
        rom[74][8] = 16'hFFB8;
        rom[74][9] = 16'hFFE1;
        rom[75][0] = 16'hFFE6;
        rom[75][1] = 16'h0022;
        rom[75][2] = 16'h0006;
        rom[75][3] = 16'hFFEA;
        rom[75][4] = 16'hFFE3;
        rom[75][5] = 16'h001D;
        rom[75][6] = 16'hFFB5;
        rom[75][7] = 16'h0001;
        rom[75][8] = 16'hFFDD;
        rom[75][9] = 16'hFFF2;
        rom[76][0] = 16'hFFD1;
        rom[76][1] = 16'hFFDC;
        rom[76][2] = 16'hFFA9;
        rom[76][3] = 16'h0003;
        rom[76][4] = 16'h002C;
        rom[76][5] = 16'h0023;
        rom[76][6] = 16'hFFE3;
        rom[76][7] = 16'hFFE3;
        rom[76][8] = 16'h0010;
        rom[76][9] = 16'h0021;
        rom[77][0] = 16'hFFED;
        rom[77][1] = 16'hFFBB;
        rom[77][2] = 16'h0042;
        rom[77][3] = 16'hFFCB;
        rom[77][4] = 16'h0032;
        rom[77][5] = 16'hFFDE;
        rom[77][6] = 16'h003E;
        rom[77][7] = 16'hFFF3;
        rom[77][8] = 16'hFFD9;
        rom[77][9] = 16'hFFFA;
        rom[78][0] = 16'h0014;
        rom[78][1] = 16'h0029;
        rom[78][2] = 16'hFFC6;
        rom[78][3] = 16'h0003;
        rom[78][4] = 16'h0009;
        rom[78][5] = 16'h0022;
        rom[78][6] = 16'hFFFD;
        rom[78][7] = 16'hFFBE;
        rom[78][8] = 16'h0006;
        rom[78][9] = 16'h0006;
        rom[79][0] = 16'hFFF8;
        rom[79][1] = 16'h001D;
        rom[79][2] = 16'hFFCF;
        rom[79][3] = 16'hFFE0;
        rom[79][4] = 16'h0015;
        rom[79][5] = 16'hFFD3;
        rom[79][6] = 16'h003E;
        rom[79][7] = 16'hFFEC;
        rom[79][8] = 16'h0006;
        rom[79][9] = 16'hFFE5;
        rom[80][0] = 16'hFFD8;
        rom[80][1] = 16'hFFFE;
        rom[80][2] = 16'h0029;
        rom[80][3] = 16'hFFE8;
        rom[80][4] = 16'hFFD1;
        rom[80][5] = 16'hFFE0;
        rom[80][6] = 16'hFFBE;
        rom[80][7] = 16'h001F;
        rom[80][8] = 16'h0027;
        rom[80][9] = 16'h0007;
        rom[81][0] = 16'hFFDC;
        rom[81][1] = 16'h0027;
        rom[81][2] = 16'hFFA7;
        rom[81][3] = 16'h002C;
        rom[81][4] = 16'hFFB7;
        rom[81][5] = 16'h0028;
        rom[81][6] = 16'hFFCA;
        rom[81][7] = 16'h0026;
        rom[81][8] = 16'hFFEB;
        rom[81][9] = 16'hFFE4;
        rom[82][0] = 16'hFFD7;
        rom[82][1] = 16'hFFE8;
        rom[82][2] = 16'hFFDA;
        rom[82][3] = 16'hFFE1;
        rom[82][4] = 16'h0016;
        rom[82][5] = 16'hFFC9;
        rom[82][6] = 16'hFFDA;
        rom[82][7] = 16'h0034;
        rom[82][8] = 16'h0031;
        rom[82][9] = 16'hFFE6;
        rom[83][0] = 16'h0027;
        rom[83][1] = 16'h0015;
        rom[83][2] = 16'h0021;
        rom[83][3] = 16'h0026;
        rom[83][4] = 16'h0003;
        rom[83][5] = 16'h002A;
        rom[83][6] = 16'h002B;
        rom[83][7] = 16'hFFDC;
        rom[83][8] = 16'h0023;
        rom[83][9] = 16'hFFDE;
        rom[84][0] = 16'hFFBC;
        rom[84][1] = 16'h0026;
        rom[84][2] = 16'hFFB8;
        rom[84][3] = 16'h0037;
        rom[84][4] = 16'hFFF4;
        rom[84][5] = 16'hFFF2;
        rom[84][6] = 16'hFFBF;
        rom[84][7] = 16'hFFF6;
        rom[84][8] = 16'hFFDB;
        rom[84][9] = 16'hFFF3;
        rom[85][0] = 16'hFFE7;
        rom[85][1] = 16'hFFC0;
        rom[85][2] = 16'hFFD3;
        rom[85][3] = 16'hFFE2;
        rom[85][4] = 16'h002A;
        rom[85][5] = 16'hFFF1;
        rom[85][6] = 16'hFFE3;
        rom[85][7] = 16'h0010;
        rom[85][8] = 16'hFFCE;
        rom[85][9] = 16'h0021;
        rom[86][0] = 16'h0009;
        rom[86][1] = 16'h0021;
        rom[86][2] = 16'h0004;
        rom[86][3] = 16'h002B;
        rom[86][4] = 16'hFFC4;
        rom[86][5] = 16'h002A;
        rom[86][6] = 16'h0017;
        rom[86][7] = 16'h0008;
        rom[86][8] = 16'hFFFB;
        rom[86][9] = 16'hFFB6;
        rom[87][0] = 16'h000C;
        rom[87][1] = 16'hFFF0;
        rom[87][2] = 16'hFFBC;
        rom[87][3] = 16'hFFD2;
        rom[87][4] = 16'h002B;
        rom[87][5] = 16'hFFD0;
        rom[87][6] = 16'h0013;
        rom[87][7] = 16'hFFC4;
        rom[87][8] = 16'h000B;
        rom[87][9] = 16'h0029;
        rom[88][0] = 16'hFFF8;
        rom[88][1] = 16'hFFE4;
        rom[88][2] = 16'h0017;
        rom[88][3] = 16'hFFBF;
        rom[88][4] = 16'h000F;
        rom[88][5] = 16'hFFE2;
        rom[88][6] = 16'h0056;
        rom[88][7] = 16'hFFE1;
        rom[88][8] = 16'hFFFA;
        rom[88][9] = 16'hFFAF;
        rom[89][0] = 16'hFFFF;
        rom[89][1] = 16'h0005;
        rom[89][2] = 16'hFFBA;
        rom[89][3] = 16'h0003;
        rom[89][4] = 16'h0029;
        rom[89][5] = 16'h0027;
        rom[89][6] = 16'h001D;
        rom[89][7] = 16'hFFBA;
        rom[89][8] = 16'hFFC9;
        rom[89][9] = 16'h002A;
        rom[90][0] = 16'hFFF0;
        rom[90][1] = 16'hFFDC;
        rom[90][2] = 16'hFFEA;
        rom[90][3] = 16'hFFEF;
        rom[90][4] = 16'h000E;
        rom[90][5] = 16'hFFD4;
        rom[90][6] = 16'h001E;
        rom[90][7] = 16'h0020;
        rom[90][8] = 16'h0027;
        rom[90][9] = 16'hFFE7;
        rom[91][0] = 16'hFFFC;
        rom[91][1] = 16'h003F;
        rom[91][2] = 16'hFFDF;
        rom[91][3] = 16'hFFE9;
        rom[91][4] = 16'h0009;
        rom[91][5] = 16'hFFE6;
        rom[91][6] = 16'hFFF9;
        rom[91][7] = 16'h0028;
        rom[91][8] = 16'h0005;
        rom[91][9] = 16'h0030;
        rom[92][0] = 16'h000F;
        rom[92][1] = 16'h000E;
        rom[92][2] = 16'hFFD8;
        rom[92][3] = 16'hFFE0;
        rom[92][4] = 16'h0020;
        rom[92][5] = 16'h0011;
        rom[92][6] = 16'hFFD9;
        rom[92][7] = 16'hFFC9;
        rom[92][8] = 16'hFFE3;
        rom[92][9] = 16'h0024;
        rom[93][0] = 16'hFFF7;
        rom[93][1] = 16'h001F;
        rom[93][2] = 16'hFFD5;
        rom[93][3] = 16'h0037;
        rom[93][4] = 16'h000B;
        rom[93][5] = 16'h0032;
        rom[93][6] = 16'hFFC9;
        rom[93][7] = 16'hFFB8;
        rom[93][8] = 16'hFFCB;
        rom[93][9] = 16'h0025;
        rom[94][0] = 16'hFFED;
        rom[94][1] = 16'hFFD9;
        rom[94][2] = 16'h002A;
        rom[94][3] = 16'h001D;
        rom[94][4] = 16'hFFDE;
        rom[94][5] = 16'hFFDD;
        rom[94][6] = 16'hFFD5;
        rom[94][7] = 16'hFFDF;
        rom[94][8] = 16'hFFFF;
        rom[94][9] = 16'hFFD5;
        rom[95][0] = 16'h0025;
        rom[95][1] = 16'hFFF3;
        rom[95][2] = 16'hFFA4;
        rom[95][3] = 16'hFFE1;
        rom[95][4] = 16'h0017;
        rom[95][5] = 16'h0033;
        rom[95][6] = 16'hFFBD;
        rom[95][7] = 16'hFFC9;
        rom[95][8] = 16'hFFC6;
        rom[95][9] = 16'h0022;
        rom[96][0] = 16'hFFDB;
        rom[96][1] = 16'h0029;
        rom[96][2] = 16'hFFDD;
        rom[96][3] = 16'h000E;
        rom[96][4] = 16'h0028;
        rom[96][5] = 16'h0031;
        rom[96][6] = 16'hFFD8;
        rom[96][7] = 16'hFFCC;
        rom[96][8] = 16'hFFEA;
        rom[96][9] = 16'h0027;
        rom[97][0] = 16'hFFE0;
        rom[97][1] = 16'h0012;
        rom[97][2] = 16'hFFC8;
        rom[97][3] = 16'hFFC4;
        rom[97][4] = 16'h001E;
        rom[97][5] = 16'h0002;
        rom[97][6] = 16'hFFE9;
        rom[97][7] = 16'h002B;
        rom[97][8] = 16'hFFD9;
        rom[97][9] = 16'hFFF6;
        rom[98][0] = 16'hFFB2;
        rom[98][1] = 16'h0027;
        rom[98][2] = 16'hFFF7;
        rom[98][3] = 16'h001D;
        rom[98][4] = 16'hFFEB;
        rom[98][5] = 16'hFFD0;
        rom[98][6] = 16'h0018;
        rom[98][7] = 16'h001C;
        rom[98][8] = 16'hFFF5;
        rom[98][9] = 16'hFFB8;
        rom[99][0] = 16'h001C;
        rom[99][1] = 16'h0028;
        rom[99][2] = 16'hFFC4;
        rom[99][3] = 16'h002C;
        rom[99][4] = 16'hFFC3;
        rom[99][5] = 16'h001D;
        rom[99][6] = 16'hFFDC;
        rom[99][7] = 16'h0023;
        rom[99][8] = 16'hFFF9;
        rom[99][9] = 16'hFFC9;
        rom[100][0] = 16'hFFBA;
        rom[100][1] = 16'h0018;
        rom[100][2] = 16'h0008;
        rom[100][3] = 16'h0005;
        rom[100][4] = 16'hFFC4;
        rom[100][5] = 16'h0014;
        rom[100][6] = 16'hFFA8;
        rom[100][7] = 16'h0028;
        rom[100][8] = 16'hFFC6;
        rom[100][9] = 16'h0004;
        rom[101][0] = 16'hFFF8;
        rom[101][1] = 16'h000A;
        rom[101][2] = 16'hFFED;
        rom[101][3] = 16'hFFCF;
        rom[101][4] = 16'h0018;
        rom[101][5] = 16'h0020;
        rom[101][6] = 16'h0014;
        rom[101][7] = 16'hFFDC;
        rom[101][8] = 16'h0027;
        rom[101][9] = 16'h0048;
        rom[102][0] = 16'hFFCE;
        rom[102][1] = 16'hFFC9;
        rom[102][2] = 16'h001D;
        rom[102][3] = 16'hFFFA;
        rom[102][4] = 16'h001C;
        rom[102][5] = 16'h0003;
        rom[102][6] = 16'hFFE4;
        rom[102][7] = 16'h003C;
        rom[102][8] = 16'hFFFF;
        rom[102][9] = 16'h0039;
        rom[103][0] = 16'h0015;
        rom[103][1] = 16'h0002;
        rom[103][2] = 16'h000B;
        rom[103][3] = 16'hFFF6;
        rom[103][4] = 16'h0031;
        rom[103][5] = 16'hFFFF;
        rom[103][6] = 16'hFFCC;
        rom[103][7] = 16'hFFCF;
        rom[103][8] = 16'hFFD9;
        rom[103][9] = 16'h003F;
        rom[104][0] = 16'hFFF1;
        rom[104][1] = 16'hFFF7;
        rom[104][2] = 16'h0008;
        rom[104][3] = 16'hFFCC;
        rom[104][4] = 16'h0036;
        rom[104][5] = 16'hFFD8;
        rom[104][6] = 16'h002C;
        rom[104][7] = 16'hFFFD;
        rom[104][8] = 16'hFFE3;
        rom[104][9] = 16'h0034;
        rom[105][0] = 16'h0066;
        rom[105][1] = 16'hFFF0;
        rom[105][2] = 16'h000D;
        rom[105][3] = 16'hFFD9;
        rom[105][4] = 16'hFFBF;
        rom[105][5] = 16'hFFCE;
        rom[105][6] = 16'hFFE5;
        rom[105][7] = 16'hFFEE;
        rom[105][8] = 16'hFFBE;
        rom[105][9] = 16'hFFF1;
        rom[106][0] = 16'hFFC2;
        rom[106][1] = 16'hFFEF;
        rom[106][2] = 16'h0009;
        rom[106][3] = 16'h0027;
        rom[106][4] = 16'h000E;
        rom[106][5] = 16'h001D;
        rom[106][6] = 16'hFFB4;
        rom[106][7] = 16'h002C;
        rom[106][8] = 16'h002A;
        rom[106][9] = 16'h0023;
        rom[107][0] = 16'hFFAF;
        rom[107][1] = 16'hFFDE;
        rom[107][2] = 16'hFFB1;
        rom[107][3] = 16'h0006;
        rom[107][4] = 16'hFFD8;
        rom[107][5] = 16'h0001;
        rom[107][6] = 16'h000B;
        rom[107][7] = 16'hFFBD;
        rom[107][8] = 16'hFFED;
        rom[107][9] = 16'hFFFD;
        rom[108][0] = 16'hFFFD;
        rom[108][1] = 16'hFFD0;
        rom[108][2] = 16'h0066;
        rom[108][3] = 16'hFFED;
        rom[108][4] = 16'h0010;
        rom[108][5] = 16'hFFD4;
        rom[108][6] = 16'h0037;
        rom[108][7] = 16'h0046;
        rom[108][8] = 16'hFFF4;
        rom[108][9] = 16'h0037;
        rom[109][0] = 16'hFFB7;
        rom[109][1] = 16'hFFEA;
        rom[109][2] = 16'hFFF8;
        rom[109][3] = 16'h0023;
        rom[109][4] = 16'h0023;
        rom[109][5] = 16'h0027;
        rom[109][6] = 16'hFFEB;
        rom[109][7] = 16'h002C;
        rom[109][8] = 16'hFFDB;
        rom[109][9] = 16'h002F;
        rom[110][0] = 16'hFFDE;
        rom[110][1] = 16'hFFE9;
        rom[110][2] = 16'hFFE5;
        rom[110][3] = 16'h0019;
        rom[110][4] = 16'h0013;
        rom[110][5] = 16'hFFF9;
        rom[110][6] = 16'hFFE0;
        rom[110][7] = 16'h001D;
        rom[110][8] = 16'h0021;
        rom[110][9] = 16'hFFE5;
        rom[111][0] = 16'hFFBA;
        rom[111][1] = 16'h0014;
        rom[111][2] = 16'hFFBA;
        rom[111][3] = 16'h001F;
        rom[111][4] = 16'hFFAF;
        rom[111][5] = 16'h0012;
        rom[111][6] = 16'hFF97;
        rom[111][7] = 16'hFFFB;
        rom[111][8] = 16'h0009;
        rom[111][9] = 16'hFFE7;
        rom[112][0] = 16'h0053;
        rom[112][1] = 16'hFFE1;
        rom[112][2] = 16'hFFFA;
        rom[112][3] = 16'hFFDE;
        rom[112][4] = 16'h0008;
        rom[112][5] = 16'hFFE9;
        rom[112][6] = 16'hFFCF;
        rom[112][7] = 16'h0028;
        rom[112][8] = 16'h0043;
        rom[112][9] = 16'hFFE9;
        rom[113][0] = 16'h0037;
        rom[113][1] = 16'hFFE5;
        rom[113][2] = 16'hFFC9;
        rom[113][3] = 16'hFFC7;
        rom[113][4] = 16'hFFC9;
        rom[113][5] = 16'hFFCE;
        rom[113][6] = 16'h0026;
        rom[113][7] = 16'hFFF9;
        rom[113][8] = 16'h0007;
        rom[113][9] = 16'hFFC7;
        rom[114][0] = 16'hFFDE;
        rom[114][1] = 16'hFFFC;
        rom[114][2] = 16'h0014;
        rom[114][3] = 16'h001D;
        rom[114][4] = 16'h001B;
        rom[114][5] = 16'hFFD5;
        rom[114][6] = 16'hFFF2;
        rom[114][7] = 16'h0024;
        rom[114][8] = 16'hFFE8;
        rom[114][9] = 16'h001D;
        rom[115][0] = 16'h003B;
        rom[115][1] = 16'h000E;
        rom[115][2] = 16'h003D;
        rom[115][3] = 16'hFFD2;
        rom[115][4] = 16'hFFCC;
        rom[115][5] = 16'hFFE2;
        rom[115][6] = 16'hFFCB;
        rom[115][7] = 16'hFFDE;
        rom[115][8] = 16'hFFCE;
        rom[115][9] = 16'hFFF7;
        rom[116][0] = 16'hFFE8;
        rom[116][1] = 16'h001C;
        rom[116][2] = 16'hFFC2;
        rom[116][3] = 16'hFFF8;
        rom[116][4] = 16'h003A;
        rom[116][5] = 16'hFFED;
        rom[116][6] = 16'hFFE1;
        rom[116][7] = 16'h0006;
        rom[116][8] = 16'hFFF8;
        rom[116][9] = 16'h0036;
        rom[117][0] = 16'h0008;
        rom[117][1] = 16'h0032;
        rom[117][2] = 16'hFFEA;
        rom[117][3] = 16'h0006;
        rom[117][4] = 16'hFFFC;
        rom[117][5] = 16'h002C;
        rom[117][6] = 16'hFFCC;
        rom[117][7] = 16'h002A;
        rom[117][8] = 16'h0026;
        rom[117][9] = 16'hFFE7;
        rom[118][0] = 16'hFFED;
        rom[118][1] = 16'hFFE0;
        rom[118][2] = 16'hFFDE;
        rom[118][3] = 16'hFFE7;
        rom[118][4] = 16'h000E;
        rom[118][5] = 16'h0012;
        rom[118][6] = 16'hFFEF;
        rom[118][7] = 16'h003B;
        rom[118][8] = 16'h0016;
        rom[118][9] = 16'hFFE2;
        rom[119][0] = 16'hFFED;
        rom[119][1] = 16'h0023;
        rom[119][2] = 16'h0001;
        rom[119][3] = 16'h002B;
        rom[119][4] = 16'hFFD1;
        rom[119][5] = 16'h002C;
        rom[119][6] = 16'hFFA6;
        rom[119][7] = 16'h0015;
        rom[119][8] = 16'hFFFC;
        rom[119][9] = 16'hFFB3;
        rom[120][0] = 16'h0032;
        rom[120][1] = 16'hFFF8;
        rom[120][2] = 16'hFFE3;
        rom[120][3] = 16'h0024;
        rom[120][4] = 16'h002E;
        rom[120][5] = 16'h0012;
        rom[120][6] = 16'h0031;
        rom[120][7] = 16'hFFD3;
        rom[120][8] = 16'hFFF2;
        rom[120][9] = 16'h001B;
        rom[121][0] = 16'hFFBC;
        rom[121][1] = 16'h0013;
        rom[121][2] = 16'hFFC2;
        rom[121][3] = 16'h0017;
        rom[121][4] = 16'hFFE1;
        rom[121][5] = 16'hFFF8;
        rom[121][6] = 16'hFFB9;
        rom[121][7] = 16'h001F;
        rom[121][8] = 16'hFFC1;
        rom[121][9] = 16'hFFB6;
        rom[122][0] = 16'hFFCD;
        rom[122][1] = 16'hFFD4;
        rom[122][2] = 16'hFFD0;
        rom[122][3] = 16'hFFD4;
        rom[122][4] = 16'h0023;
        rom[122][5] = 16'hFFFD;
        rom[122][6] = 16'h0032;
        rom[122][7] = 16'hFFC2;
        rom[122][8] = 16'hFFE4;
        rom[122][9] = 16'h0027;
        rom[123][0] = 16'h0006;
        rom[123][1] = 16'h002F;
        rom[123][2] = 16'hFFC5;
        rom[123][3] = 16'h0000;
        rom[123][4] = 16'h0022;
        rom[123][5] = 16'h001A;
        rom[123][6] = 16'hFFAE;
        rom[123][7] = 16'hFFFD;
        rom[123][8] = 16'hFFA7;
        rom[123][9] = 16'h003C;
        rom[124][0] = 16'hFFF8;
        rom[124][1] = 16'h0027;
        rom[124][2] = 16'hFFD6;
        rom[124][3] = 16'hFFFD;
        rom[124][4] = 16'h0027;
        rom[124][5] = 16'h001D;
        rom[124][6] = 16'hFFEB;
        rom[124][7] = 16'hFFD4;
        rom[124][8] = 16'hFFE7;
        rom[124][9] = 16'h002F;
        rom[125][0] = 16'hFFE0;
        rom[125][1] = 16'hFFF2;
        rom[125][2] = 16'hFFA2;
        rom[125][3] = 16'hFFD2;
        rom[125][4] = 16'h002E;
        rom[125][5] = 16'hFFEF;
        rom[125][6] = 16'h002C;
        rom[125][7] = 16'h0004;
        rom[125][8] = 16'h0017;
        rom[125][9] = 16'h0025;
        rom[126][0] = 16'hFFD6;
        rom[126][1] = 16'h000B;
        rom[126][2] = 16'h0026;
        rom[126][3] = 16'hFFE8;
        rom[126][4] = 16'h0002;
        rom[126][5] = 16'hFFD5;
        rom[126][6] = 16'hFFFC;
        rom[126][7] = 16'h004F;
        rom[126][8] = 16'hFFDD;
        rom[126][9] = 16'h0027;
        rom[127][0] = 16'h0020;
        rom[127][1] = 16'h0015;
        rom[127][2] = 16'hFFDE;
        rom[127][3] = 16'h0000;
        rom[127][4] = 16'h0006;
        rom[127][5] = 16'hFFD4;
        rom[127][6] = 16'h0023;
        rom[127][7] = 16'hFFDD;
        rom[127][8] = 16'h0001;
        rom[127][9] = 16'h002A;
    end

    always @(*) begin
        data_out = rom[addr][index];
    end
endmodule
