// Q8.8 Fixed-Point ROM: rom_layer0_biases
module rom_layer0_biases (
    input [7:0] addr,
    output reg signed [15:0] data_out
);

    reg signed [15:0] rom [0:255];

    initial begin
        rom[0] = 16'hFF87;
        rom[1] = 16'hFFA4;
        rom[2] = 16'hFF7B;
        rom[3] = 16'hFF9A;
        rom[4] = 16'hFFCB;
        rom[5] = 16'hFF80;
        rom[6] = 16'hFF63;
        rom[7] = 16'hFF7E;
        rom[8] = 16'hFF76;
        rom[9] = 16'hFFA6;
        rom[10] = 16'hFF7D;
        rom[11] = 16'hFF91;
        rom[12] = 16'hFF55;
        rom[13] = 16'hFF5E;
        rom[14] = 16'hFF95;
        rom[15] = 16'hFF8C;
        rom[16] = 16'hFF96;
        rom[17] = 16'hFF66;
        rom[18] = 16'hFF44;
        rom[19] = 16'hFF52;
        rom[20] = 16'hFF37;
        rom[21] = 16'hFF6F;
        rom[22] = 16'hFF78;
        rom[23] = 16'hFF66;
        rom[24] = 16'hFF68;
        rom[25] = 16'hFF66;
        rom[26] = 16'hFF43;
        rom[27] = 16'hFF7E;
        rom[28] = 16'hFF95;
        rom[29] = 16'hFF4D;
        rom[30] = 16'hFF93;
        rom[31] = 16'hFF89;
        rom[32] = 16'hFF8E;
        rom[33] = 16'hFF7B;
        rom[34] = 16'hFF7B;
        rom[35] = 16'hFF96;
        rom[36] = 16'hFF29;
        rom[37] = 16'hFF59;
        rom[38] = 16'hFF89;
        rom[39] = 16'hFFA0;
        rom[40] = 16'hFF96;
        rom[41] = 16'hFF61;
        rom[42] = 16'hFF63;
        rom[43] = 16'hFF48;
        rom[44] = 16'hFFC1;
        rom[45] = 16'hFF95;
        rom[46] = 16'hFF9B;
        rom[47] = 16'hFF52;
        rom[48] = 16'hFFD0;
        rom[49] = 16'hFF89;
        rom[50] = 16'hFF71;
        rom[51] = 16'hFF66;
        rom[52] = 16'hFF55;
        rom[53] = 16'hFF74;
        rom[54] = 16'hFF8F;
        rom[55] = 16'hFF65;
        rom[56] = 16'hFF79;
        rom[57] = 16'hFF8F;
        rom[58] = 16'hFF72;
        rom[59] = 16'hFF61;
        rom[60] = 16'hFF71;
        rom[61] = 16'hFF93;
        rom[62] = 16'hFF74;
        rom[63] = 16'hFF55;
        rom[64] = 16'hFF80;
        rom[65] = 16'hFFA2;
        rom[66] = 16'hFF44;
        rom[67] = 16'hFF82;
        rom[68] = 16'hFF6F;
        rom[69] = 16'hFF6D;
        rom[70] = 16'hFF8C;
        rom[71] = 16'hFF76;
        rom[72] = 16'hFF83;
        rom[73] = 16'hFF41;
        rom[74] = 16'hFF95;
        rom[75] = 16'hFF7E;
        rom[76] = 16'hFF9B;
        rom[77] = 16'hFF2B;
        rom[78] = 16'hFFA6;
        rom[79] = 16'hFF6C;
        rom[80] = 16'hFF5E;
        rom[81] = 16'hFF82;
        rom[82] = 16'hFF63;
        rom[83] = 16'hFF55;
        rom[84] = 16'hFFA2;
        rom[85] = 16'hFF8A;
        rom[86] = 16'hFF48;
        rom[87] = 16'hFF8A;
        rom[88] = 16'hFF72;
        rom[89] = 16'hFF74;
        rom[90] = 16'hFF6F;
        rom[91] = 16'hFF82;
        rom[92] = 16'hFF8E;
        rom[93] = 16'hFF8F;
        rom[94] = 16'hFF8E;
        rom[95] = 16'hFF6C;
        rom[96] = 16'hFF46;
        rom[97] = 16'hFF4B;
        rom[98] = 16'hFF4F;
        rom[99] = 16'hFFB2;
        rom[100] = 16'hFF27;
        rom[101] = 16'hFF54;
        rom[102] = 16'hFF79;
        rom[103] = 16'hFF79;
        rom[104] = 16'hFFAC;
        rom[105] = 16'hFF80;
        rom[106] = 16'hFF8E;
        rom[107] = 16'hFF80;
        rom[108] = 16'hFF6D;
        rom[109] = 16'hFF66;
        rom[110] = 16'hFF5E;
        rom[111] = 16'hFFA2;
        rom[112] = 16'hFF72;
        rom[113] = 16'hFF93;
        rom[114] = 16'hFF8A;
        rom[115] = 16'hFF66;
        rom[116] = 16'hFF87;
        rom[117] = 16'hFF71;
        rom[118] = 16'hFFA7;
        rom[119] = 16'hFF9F;
        rom[120] = 16'hFF96;
        rom[121] = 16'hFF6F;
        rom[122] = 16'hFF6D;
        rom[123] = 16'hFF85;
        rom[124] = 16'hFF96;
        rom[125] = 16'hFF9D;
        rom[126] = 16'hFF82;
        rom[127] = 16'hFF6A;
        rom[128] = 16'hFF7D;
        rom[129] = 16'hFF6A;
        rom[130] = 16'hFF48;
        rom[131] = 16'hFF4F;
        rom[132] = 16'hFF4F;
        rom[133] = 16'hFF9A;
        rom[134] = 16'hFF7D;
        rom[135] = 16'hFF60;
        rom[136] = 16'hFF95;
        rom[137] = 16'hFF63;
        rom[138] = 16'hFF85;
        rom[139] = 16'hFF89;
        rom[140] = 16'hFF41;
        rom[141] = 16'hFF6F;
        rom[142] = 16'hFF4B;
        rom[143] = 16'hFF7B;
        rom[144] = 16'hFF74;
        rom[145] = 16'hFF49;
        rom[146] = 16'hFF59;
        rom[147] = 16'hFF7E;
        rom[148] = 16'hFF66;
        rom[149] = 16'hFF6C;
        rom[150] = 16'hFF8E;
        rom[151] = 16'hFF72;
        rom[152] = 16'hFF44;
        rom[153] = 16'hFF3F;
        rom[154] = 16'hFF79;
        rom[155] = 16'hFF5B;
        rom[156] = 16'hFF74;
        rom[157] = 16'hFF6C;
        rom[158] = 16'hFF74;
        rom[159] = 16'hFF65;
        rom[160] = 16'hFF95;
        rom[161] = 16'hFF76;
        rom[162] = 16'hFF8A;
        rom[163] = 16'hFF89;
        rom[164] = 16'hFF85;
        rom[165] = 16'hFF6C;
        rom[166] = 16'hFF7B;
        rom[167] = 16'hFF8A;
        rom[168] = 16'hFF4F;
        rom[169] = 16'hFF8C;
        rom[170] = 16'hFF57;
        rom[171] = 16'hFFBC;
        rom[172] = 16'hFFA9;
        rom[173] = 16'hFF7D;
        rom[174] = 16'hFFB2;
        rom[175] = 16'hFF95;
        rom[176] = 16'hFF7B;
        rom[177] = 16'hFF68;
        rom[178] = 16'hFF55;
        rom[179] = 16'hFF71;
        rom[180] = 16'hFF7E;
        rom[181] = 16'hFF63;
        rom[182] = 16'hFF55;
        rom[183] = 16'hFF8A;
        rom[184] = 16'hFF50;
        rom[185] = 16'hFF44;
        rom[186] = 16'hFF44;
        rom[187] = 16'hFF63;
        rom[188] = 16'hFFA0;
        rom[189] = 16'hFF3E;
        rom[190] = 16'hFF49;
        rom[191] = 16'hFF7B;
        rom[192] = 16'hFF8C;
        rom[193] = 16'hFF80;
        rom[194] = 16'hFF61;
        rom[195] = 16'hFFB3;
        rom[196] = 16'hFF57;
        rom[197] = 16'hFF68;
        rom[198] = 16'hFF8A;
        rom[199] = 16'hFF8C;
        rom[200] = 16'hFF71;
        rom[201] = 16'hFF72;
        rom[202] = 16'hFF4F;
        rom[203] = 16'hFF8A;
        rom[204] = 16'hFF2C;
        rom[205] = 16'hFF8F;
        rom[206] = 16'hFF80;
        rom[207] = 16'hFF83;
        rom[208] = 16'hFF82;
        rom[209] = 16'hFF60;
        rom[210] = 16'hFFB3;
        rom[211] = 16'hFF87;
        rom[212] = 16'hFF37;
        rom[213] = 16'hFFA4;
        rom[214] = 16'hFF68;
        rom[215] = 16'hFF71;
        rom[216] = 16'hFF82;
        rom[217] = 16'hFF50;
        rom[218] = 16'hFF6D;
        rom[219] = 16'hFF87;
        rom[220] = 16'hFF7D;
        rom[221] = 16'hFF50;
        rom[222] = 16'hFF3C;
        rom[223] = 16'hFF80;
        rom[224] = 16'hFF7B;
        rom[225] = 16'hFF78;
        rom[226] = 16'hFF95;
        rom[227] = 16'hFF87;
        rom[228] = 16'hFF7E;
        rom[229] = 16'hFF83;
        rom[230] = 16'hFF33;
        rom[231] = 16'hFF57;
        rom[232] = 16'hFF7B;
        rom[233] = 16'hFF8E;
        rom[234] = 16'hFF89;
        rom[235] = 16'hFF66;
        rom[236] = 16'hFF9D;
        rom[237] = 16'hFF9D;
        rom[238] = 16'hFF8A;
        rom[239] = 16'hFF78;
        rom[240] = 16'hFF9D;
        rom[241] = 16'hFF98;
        rom[242] = 16'hFF6C;
        rom[243] = 16'hFF8E;
        rom[244] = 16'hFF85;
        rom[245] = 16'hFF72;
        rom[246] = 16'hFF87;
        rom[247] = 16'hFF78;
        rom[248] = 16'hFF82;
        rom[249] = 16'hFF46;
        rom[250] = 16'hFF87;
        rom[251] = 16'hFF89;
        rom[252] = 16'hFF78;
        rom[253] = 16'hFF89;
        rom[254] = 16'hFF6C;
        rom[255] = 16'hFF68;
    end

    always @(*) begin
        data_out = rom[addr];
    end
endmodule
